##
## LEF for PtnCells ;
## created by Innovus v20.10-p004_1 on Wed Dec 29 19:58:46 2021
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO rest_top
  CLASS BLOCK ;
  SIZE 1926.480000 BY 2595.220000 ;
  FOREIGN rest_top 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1939 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.614 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 94.408 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.9096 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 26.496 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.917 LAYER met4  ;
    ANTENNAMAXAREACAR 37.7413 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 195.563 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.992488 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 3.730000 0.000000 3.870000 0.490000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4703 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.1255 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 12.2077 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 59.8263 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1.930000 0.000000 2.070000 0.485000 ;
    END
  END wb_rst_i
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.730000 0.000000 405.870000 0.490000 ;
    END
  END wbs_stb_i
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.430000 0.000000 136.570000 0.490000 ;
    END
  END wbs_cyc_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.630000 0.000000 409.770000 0.490000 ;
    END
  END wbs_we_i
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.830000 0.000000 401.970000 0.490000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.930000 0.000000 398.070000 0.490000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.030000 0.000000 394.170000 0.490000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.130000 0.000000 390.270000 0.490000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.330000 0.000000 261.470000 0.490000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.330000 0.000000 257.470000 0.490000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.430000 0.000000 253.570000 0.490000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.630000 0.000000 249.770000 0.490000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.730000 0.000000 245.870000 0.490000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.830000 0.000000 241.970000 0.490000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.930000 0.000000 238.070000 0.490000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.030000 0.000000 234.170000 0.490000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.030000 0.000000 230.170000 0.490000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.130000 0.000000 226.270000 0.490000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.230000 0.000000 222.370000 0.490000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.430000 0.000000 218.570000 0.490000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.530000 0.000000 214.670000 0.490000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.630000 0.000000 210.770000 0.490000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.630000 0.000000 206.770000 0.490000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.730000 0.000000 202.870000 0.490000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.830000 0.000000 198.970000 0.490000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.930000 0.000000 195.070000 0.490000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.030000 0.000000 191.170000 0.490000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.130000 0.000000 187.270000 0.490000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.330000 0.000000 183.470000 0.490000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.330000 0.000000 179.470000 0.490000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.430000 0.000000 175.570000 0.490000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.530000 0.000000 171.670000 0.490000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.630000 0.000000 167.770000 0.490000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.730000 0.000000 163.870000 0.490000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.830000 0.000000 159.970000 0.490000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.930000 0.000000 156.070000 0.490000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.930000 0.000000 152.070000 0.490000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.130000 0.000000 148.270000 0.490000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.230000 0.000000 144.370000 0.490000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.330000 0.000000 140.470000 0.490000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.530000 0.000000 132.670000 0.490000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.630000 0.000000 128.770000 0.490000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.730000 0.000000 124.870000 0.490000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.830000 0.000000 120.970000 0.490000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930000 0.000000 117.070000 0.490000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.030000 0.000000 113.170000 0.490000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.130000 0.000000 109.270000 0.490000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.230000 0.000000 105.370000 0.490000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.230000 0.000000 101.370000 0.490000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.330000 0.000000 97.470000 0.490000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.430000 0.000000 93.570000 0.490000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.530000 0.000000 89.670000 0.490000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.630000 0.000000 85.770000 0.490000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.730000 0.000000 81.870000 0.490000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830000 0.000000 77.970000 0.490000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.930000 0.000000 74.070000 0.490000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.030000 0.000000 70.170000 0.490000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.130000 0.000000 66.270000 0.490000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.330000 0.000000 62.470000 0.490000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.430000 0.000000 58.570000 0.490000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.530000 0.000000 54.670000 0.490000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.530000 0.000000 50.670000 0.490000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.630000 0.000000 46.770000 0.490000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.730000 0.000000 42.870000 0.490000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.830000 0.000000 38.970000 0.490000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.930000 0.000000 35.070000 0.490000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.030000 0.000000 31.170000 0.490000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.130000 0.000000 27.270000 0.490000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.130000 0.000000 23.270000 0.490000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.230000 0.000000 19.370000 0.490000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.330000 0.000000 15.470000 0.490000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.430000 0.000000 11.570000 0.490000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_ack_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5718 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.633 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 7.530000 0.000000 7.670000 0.490000 ;
    END
  END wbs_ack_o
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9322 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.553 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 386.130000 0.000000 386.270000 0.490000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9098 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.441 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 382.230000 0.000000 382.370000 0.490000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.879 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.287 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 378.330000 0.000000 378.470000 0.490000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8958 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.371 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 374.430000 0.000000 374.570000 0.490000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 370.630000 0.000000 370.770000 0.490000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9336 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.56 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 366.730000 0.000000 366.870000 0.490000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 362.830000 0.000000 362.970000 0.490000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9364 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.574 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 358.930000 0.000000 359.070000 0.490000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 355.030000 0.000000 355.170000 0.490000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8734 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.259 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 351.130000 0.000000 351.270000 0.490000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 347.230000 0.000000 347.370000 0.490000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 343.330000 0.000000 343.470000 0.490000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 339.430000 0.000000 339.570000 0.490000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9308 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.546 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 335.430000 0.000000 335.570000 0.490000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 331.530000 0.000000 331.670000 0.490000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9336 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.56 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 327.630000 0.000000 327.770000 0.490000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9098 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.441 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 323.730000 0.000000 323.870000 0.490000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 319.830000 0.000000 319.970000 0.490000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 315.930000 0.000000 316.070000 0.490000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9392 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.588 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 312.030000 0.000000 312.170000 0.490000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 308.130000 0.000000 308.270000 0.490000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9392 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.588 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 304.230000 0.000000 304.370000 0.490000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 300.330000 0.000000 300.470000 0.490000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8762 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.273 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 296.430000 0.000000 296.570000 0.490000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 292.530000 0.000000 292.670000 0.490000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 288.730000 0.000000 288.870000 0.490000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 284.730000 0.000000 284.870000 0.490000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9308 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.546 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 280.830000 0.000000 280.970000 0.490000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9154 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.469 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 276.930000 0.000000 277.070000 0.490000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 273.030000 0.000000 273.170000 0.490000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8902 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 269.130000 0.000000 269.270000 0.490000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9252 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.518 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 265.230000 0.000000 265.370000 0.490000 ;
    END
  END wbs_dat_o[0]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 909.230000 0.000000 909.370000 0.490000 ;
    END
  END la_data_in[127]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 905.330000 0.000000 905.470000 0.490000 ;
    END
  END la_data_in[126]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.430000 0.000000 901.570000 0.490000 ;
    END
  END la_data_in[125]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 897.530000 0.000000 897.670000 0.490000 ;
    END
  END la_data_in[124]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 893.630000 0.000000 893.770000 0.490000 ;
    END
  END la_data_in[123]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.730000 0.000000 889.870000 0.490000 ;
    END
  END la_data_in[122]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 885.830000 0.000000 885.970000 0.490000 ;
    END
  END la_data_in[121]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 881.830000 0.000000 881.970000 0.490000 ;
    END
  END la_data_in[120]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.930000 0.000000 878.070000 0.490000 ;
    END
  END la_data_in[119]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 874.030000 0.000000 874.170000 0.490000 ;
    END
  END la_data_in[118]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 870.130000 0.000000 870.270000 0.490000 ;
    END
  END la_data_in[117]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 866.330000 0.000000 866.470000 0.490000 ;
    END
  END la_data_in[116]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 862.530000 0.000000 862.670000 0.490000 ;
    END
  END la_data_in[115]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 858.630000 0.000000 858.770000 0.490000 ;
    END
  END la_data_in[114]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 854.630000 0.000000 854.770000 0.490000 ;
    END
  END la_data_in[113]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.730000 0.000000 850.870000 0.490000 ;
    END
  END la_data_in[112]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.830000 0.000000 846.970000 0.490000 ;
    END
  END la_data_in[111]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 842.930000 0.000000 843.070000 0.490000 ;
    END
  END la_data_in[110]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 839.030000 0.000000 839.170000 0.490000 ;
    END
  END la_data_in[109]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.130000 0.000000 835.270000 0.490000 ;
    END
  END la_data_in[108]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 831.130000 0.000000 831.270000 0.490000 ;
    END
  END la_data_in[107]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 827.230000 0.000000 827.370000 0.490000 ;
    END
  END la_data_in[106]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 823.330000 0.000000 823.470000 0.490000 ;
    END
  END la_data_in[105]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 819.430000 0.000000 819.570000 0.490000 ;
    END
  END la_data_in[104]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.530000 0.000000 815.670000 0.490000 ;
    END
  END la_data_in[103]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.630000 0.000000 811.770000 0.490000 ;
    END
  END la_data_in[102]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 807.730000 0.000000 807.870000 0.490000 ;
    END
  END la_data_in[101]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 803.830000 0.000000 803.970000 0.490000 ;
    END
  END la_data_in[100]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 799.930000 0.000000 800.070000 0.490000 ;
    END
  END la_data_in[99]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 796.030000 0.000000 796.170000 0.490000 ;
    END
  END la_data_in[98]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.230000 0.000000 792.370000 0.490000 ;
    END
  END la_data_in[97]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.330000 0.000000 788.470000 0.490000 ;
    END
  END la_data_in[96]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.430000 0.000000 784.570000 0.490000 ;
    END
  END la_data_in[95]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 780.530000 0.000000 780.670000 0.490000 ;
    END
  END la_data_in[94]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.530000 0.000000 776.670000 0.490000 ;
    END
  END la_data_in[93]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.630000 0.000000 772.770000 0.490000 ;
    END
  END la_data_in[92]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 768.730000 0.000000 768.870000 0.490000 ;
    END
  END la_data_in[91]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.830000 0.000000 764.970000 0.490000 ;
    END
  END la_data_in[90]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.930000 0.000000 761.070000 0.490000 ;
    END
  END la_data_in[89]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 757.030000 0.000000 757.170000 0.490000 ;
    END
  END la_data_in[88]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.030000 0.000000 753.170000 0.490000 ;
    END
  END la_data_in[87]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.130000 0.000000 749.270000 0.490000 ;
    END
  END la_data_in[86]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.230000 0.000000 745.370000 0.490000 ;
    END
  END la_data_in[85]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.430000 0.000000 741.570000 0.490000 ;
    END
  END la_data_in[84]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.530000 0.000000 737.670000 0.490000 ;
    END
  END la_data_in[83]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.630000 0.000000 733.770000 0.490000 ;
    END
  END la_data_in[82]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.730000 0.000000 729.870000 0.490000 ;
    END
  END la_data_in[81]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.730000 0.000000 725.870000 0.490000 ;
    END
  END la_data_in[80]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.930000 0.000000 722.070000 0.490000 ;
    END
  END la_data_in[79]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.030000 0.000000 718.170000 0.490000 ;
    END
  END la_data_in[78]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.130000 0.000000 714.270000 0.490000 ;
    END
  END la_data_in[77]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.230000 0.000000 710.370000 0.490000 ;
    END
  END la_data_in[76]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.330000 0.000000 706.470000 0.490000 ;
    END
  END la_data_in[75]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.430000 0.000000 702.570000 0.490000 ;
    END
  END la_data_in[74]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.430000 0.000000 698.570000 0.490000 ;
    END
  END la_data_in[73]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.530000 0.000000 694.670000 0.490000 ;
    END
  END la_data_in[72]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.630000 0.000000 690.770000 0.490000 ;
    END
  END la_data_in[71]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.730000 0.000000 686.870000 0.490000 ;
    END
  END la_data_in[70]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.830000 0.000000 682.970000 0.490000 ;
    END
  END la_data_in[69]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.930000 0.000000 679.070000 0.490000 ;
    END
  END la_data_in[68]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 675.030000 0.000000 675.170000 0.490000 ;
    END
  END la_data_in[67]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 671.130000 0.000000 671.270000 0.490000 ;
    END
  END la_data_in[66]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.230000 0.000000 667.370000 0.490000 ;
    END
  END la_data_in[65]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.330000 0.000000 663.470000 0.490000 ;
    END
  END la_data_in[64]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 659.430000 0.000000 659.570000 0.490000 ;
    END
  END la_data_in[63]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 655.530000 0.000000 655.670000 0.490000 ;
    END
  END la_data_in[62]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 651.630000 0.000000 651.770000 0.490000 ;
    END
  END la_data_in[61]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.730000 0.000000 647.870000 0.490000 ;
    END
  END la_data_in[60]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.830000 0.000000 643.970000 0.490000 ;
    END
  END la_data_in[59]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.930000 0.000000 640.070000 0.490000 ;
    END
  END la_data_in[58]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 636.030000 0.000000 636.170000 0.490000 ;
    END
  END la_data_in[57]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.130000 0.000000 632.270000 0.490000 ;
    END
  END la_data_in[56]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.230000 0.000000 628.370000 0.490000 ;
    END
  END la_data_in[55]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.330000 0.000000 624.470000 0.490000 ;
    END
  END la_data_in[54]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.430000 0.000000 620.570000 0.490000 ;
    END
  END la_data_in[53]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.530000 0.000000 616.670000 0.490000 ;
    END
  END la_data_in[52]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.630000 0.000000 612.770000 0.490000 ;
    END
  END la_data_in[51]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.730000 0.000000 608.870000 0.490000 ;
    END
  END la_data_in[50]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.830000 0.000000 604.970000 0.490000 ;
    END
  END la_data_in[49]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 600.930000 0.000000 601.070000 0.490000 ;
    END
  END la_data_in[48]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 596.930000 0.000000 597.070000 0.490000 ;
    END
  END la_data_in[47]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.030000 0.000000 593.170000 0.490000 ;
    END
  END la_data_in[46]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.130000 0.000000 589.270000 0.490000 ;
    END
  END la_data_in[45]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.230000 0.000000 585.370000 0.490000 ;
    END
  END la_data_in[44]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.330000 0.000000 581.470000 0.490000 ;
    END
  END la_data_in[43]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.530000 0.000000 577.670000 0.490000 ;
    END
  END la_data_in[42]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.630000 0.000000 573.770000 0.490000 ;
    END
  END la_data_in[41]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.630000 0.000000 569.770000 0.490000 ;
    END
  END la_data_in[40]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.730000 0.000000 565.870000 0.490000 ;
    END
  END la_data_in[39]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.830000 0.000000 561.970000 0.490000 ;
    END
  END la_data_in[38]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.930000 0.000000 558.070000 0.490000 ;
    END
  END la_data_in[37]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 554.130000 0.000000 554.270000 0.490000 ;
    END
  END la_data_in[36]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.230000 0.000000 550.370000 0.490000 ;
    END
  END la_data_in[35]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.330000 0.000000 546.470000 0.490000 ;
    END
  END la_data_in[34]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.330000 0.000000 542.470000 0.490000 ;
    END
  END la_data_in[33]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.430000 0.000000 538.570000 0.490000 ;
    END
  END la_data_in[32]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.530000 0.000000 534.670000 0.490000 ;
    END
  END la_data_in[31]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.630000 0.000000 530.770000 0.490000 ;
    END
  END la_data_in[30]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.730000 0.000000 526.870000 0.490000 ;
    END
  END la_data_in[29]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.830000 0.000000 522.970000 0.490000 ;
    END
  END la_data_in[28]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.830000 0.000000 518.970000 0.490000 ;
    END
  END la_data_in[27]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.930000 0.000000 515.070000 0.490000 ;
    END
  END la_data_in[26]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.030000 0.000000 511.170000 0.490000 ;
    END
  END la_data_in[25]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.230000 0.000000 507.370000 0.490000 ;
    END
  END la_data_in[24]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.330000 0.000000 503.470000 0.490000 ;
    END
  END la_data_in[23]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.430000 0.000000 499.570000 0.490000 ;
    END
  END la_data_in[22]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.530000 0.000000 495.670000 0.490000 ;
    END
  END la_data_in[21]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.630000 0.000000 491.770000 0.490000 ;
    END
  END la_data_in[20]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.730000 0.000000 487.870000 0.490000 ;
    END
  END la_data_in[19]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.830000 0.000000 483.970000 0.490000 ;
    END
  END la_data_in[18]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.930000 0.000000 480.070000 0.490000 ;
    END
  END la_data_in[17]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.030000 0.000000 476.170000 0.490000 ;
    END
  END la_data_in[16]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.635 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.067 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 35.2861 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 166.187 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 472.130000 0.000000 472.270000 0.490000 ;
    END
  END la_data_in[15]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9283 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.5335 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 35.6694 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 168.103 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 468.230000 0.000000 468.370000 0.490000 ;
    END
  END la_data_in[14]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6924 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.354 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 34.2321 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 155.345 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 464.230000 0.000000 464.370000 0.490000 ;
    END
  END la_data_in[13]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3718 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.751 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 14.9154 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 72.6081 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 460.330000 0.000000 460.470000 0.490000 ;
    END
  END la_data_in[12]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4054 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.919 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 14.7909 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 71.9859 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 456.430000 0.000000 456.570000 0.490000 ;
    END
  END la_data_in[11]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3059 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.5008 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.808 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 61.5612 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 313.923 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 452.530000 0.000000 452.670000 0.490000 ;
    END
  END la_data_in[10]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3956 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.87 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 30.9639 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 144.575 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 448.630000 0.000000 448.770000 0.490000 ;
    END
  END la_data_in[9]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.921 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.379 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 25.0372 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 121.889 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 444.730000 0.000000 444.870000 0.490000 ;
    END
  END la_data_in[8]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7918 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.851 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 17.2661 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 80.5111 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 440.730000 0.000000 440.870000 0.490000 ;
    END
  END la_data_in[7]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7764 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.774 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 16.1665 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 78.7455 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 436.930000 0.000000 437.070000 0.490000 ;
    END
  END la_data_in[6]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.553 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.657 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 32.7774 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 160.253 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 433.130000 0.000000 433.270000 0.490000 ;
    END
  END la_data_in[5]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.2054 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.919 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 34.6267 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 167.618 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 429.230000 0.000000 429.370000 0.490000 ;
    END
  END la_data_in[4]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3634 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.709 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 17.1982 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 81.1333 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 425.330000 0.000000 425.470000 0.490000 ;
    END
  END la_data_in[3]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.425 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.017 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 14.8701 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 72.3818 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 421.430000 0.000000 421.570000 0.490000 ;
    END
  END la_data_in[2]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.867 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.227 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 24.4788 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 116.879 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 417.530000 0.000000 417.670000 0.490000 ;
    END
  END la_data_in[1]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.103 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.407 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 13.7877 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 65.5455 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 413.530000 0.000000 413.670000 0.490000 ;
    END
  END la_data_in[0]
  PIN la_data_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9014 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.399 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1408.930000 0.000000 1409.070000 0.490000 ;
    END
  END la_data_out[127]
  PIN la_data_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9322 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.553 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1405.030000 0.000000 1405.170000 0.490000 ;
    END
  END la_data_out[126]
  PIN la_data_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8958 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.371 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1401.030000 0.000000 1401.170000 0.490000 ;
    END
  END la_data_out[125]
  PIN la_data_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.879 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.287 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1397.130000 0.000000 1397.270000 0.490000 ;
    END
  END la_data_out[124]
  PIN la_data_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9098 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.441 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1393.230000 0.000000 1393.370000 0.490000 ;
    END
  END la_data_out[123]
  PIN la_data_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9322 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.553 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1389.330000 0.000000 1389.470000 0.490000 ;
    END
  END la_data_out[122]
  PIN la_data_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9014 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.399 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1385.430000 0.000000 1385.570000 0.490000 ;
    END
  END la_data_out[121]
  PIN la_data_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.935 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.567 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1381.530000 0.000000 1381.670000 0.490000 ;
    END
  END la_data_out[120]
  PIN la_data_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8902 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1377.530000 0.000000 1377.670000 0.490000 ;
    END
  END la_data_out[119]
  PIN la_data_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9238 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.511 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1373.630000 0.000000 1373.770000 0.490000 ;
    END
  END la_data_out[118]
  PIN la_data_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.907 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.427 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1369.830000 0.000000 1369.970000 0.490000 ;
    END
  END la_data_out[117]
  PIN la_data_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8762 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.273 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1365.930000 0.000000 1366.070000 0.490000 ;
    END
  END la_data_out[116]
  PIN la_data_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8986 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.385 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1362.030000 0.000000 1362.170000 0.490000 ;
    END
  END la_data_out[115]
  PIN la_data_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.879 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.287 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1358.130000 0.000000 1358.270000 0.490000 ;
    END
  END la_data_out[114]
  PIN la_data_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9126 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.455 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1354.230000 0.000000 1354.370000 0.490000 ;
    END
  END la_data_out[113]
  PIN la_data_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8818 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.301 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1350.330000 0.000000 1350.470000 0.490000 ;
    END
  END la_data_out[112]
  PIN la_data_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9154 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.469 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1346.430000 0.000000 1346.570000 0.490000 ;
    END
  END la_data_out[111]
  PIN la_data_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8846 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.315 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1342.530000 0.000000 1342.670000 0.490000 ;
    END
  END la_data_out[110]
  PIN la_data_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9182 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.483 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1338.630000 0.000000 1338.770000 0.490000 ;
    END
  END la_data_out[109]
  PIN la_data_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8874 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.329 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1334.730000 0.000000 1334.870000 0.490000 ;
    END
  END la_data_out[108]
  PIN la_data_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.921 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.497 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1330.830000 0.000000 1330.970000 0.490000 ;
    END
  END la_data_out[107]
  PIN la_data_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9196 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.49 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1326.930000 0.000000 1327.070000 0.490000 ;
    END
  END la_data_out[106]
  PIN la_data_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1322.930000 0.000000 1323.070000 0.490000 ;
    END
  END la_data_out[105]
  PIN la_data_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9336 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.56 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1319.030000 0.000000 1319.170000 0.490000 ;
    END
  END la_data_out[104]
  PIN la_data_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1315.130000 0.000000 1315.270000 0.490000 ;
    END
  END la_data_out[103]
  PIN la_data_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9308 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.546 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1311.230000 0.000000 1311.370000 0.490000 ;
    END
  END la_data_out[102]
  PIN la_data_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1307.330000 0.000000 1307.470000 0.490000 ;
    END
  END la_data_out[101]
  PIN la_data_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8846 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.315 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1303.430000 0.000000 1303.570000 0.490000 ;
    END
  END la_data_out[100]
  PIN la_data_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1299.530000 0.000000 1299.670000 0.490000 ;
    END
  END la_data_out[99]
  PIN la_data_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1295.730000 0.000000 1295.870000 0.490000 ;
    END
  END la_data_out[98]
  PIN la_data_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9392 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.588 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1291.830000 0.000000 1291.970000 0.490000 ;
    END
  END la_data_out[97]
  PIN la_data_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.413 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1287.930000 0.000000 1288.070000 0.490000 ;
    END
  END la_data_out[96]
  PIN la_data_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9392 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.588 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1284.030000 0.000000 1284.170000 0.490000 ;
    END
  END la_data_out[95]
  PIN la_data_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1280.130000 0.000000 1280.270000 0.490000 ;
    END
  END la_data_out[94]
  PIN la_data_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9364 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.574 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1276.230000 0.000000 1276.370000 0.490000 ;
    END
  END la_data_out[93]
  PIN la_data_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1272.230000 0.000000 1272.370000 0.490000 ;
    END
  END la_data_out[92]
  PIN la_data_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9336 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.56 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1268.330000 0.000000 1268.470000 0.490000 ;
    END
  END la_data_out[91]
  PIN la_data_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1264.430000 0.000000 1264.570000 0.490000 ;
    END
  END la_data_out[90]
  PIN la_data_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9364 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.574 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1260.530000 0.000000 1260.670000 0.490000 ;
    END
  END la_data_out[89]
  PIN la_data_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1256.630000 0.000000 1256.770000 0.490000 ;
    END
  END la_data_out[88]
  PIN la_data_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1252.730000 0.000000 1252.870000 0.490000 ;
    END
  END la_data_out[87]
  PIN la_data_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.413 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1248.830000 0.000000 1248.970000 0.490000 ;
    END
  END la_data_out[86]
  PIN la_data_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1244.830000 0.000000 1244.970000 0.490000 ;
    END
  END la_data_out[85]
  PIN la_data_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9154 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.469 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1240.930000 0.000000 1241.070000 0.490000 ;
    END
  END la_data_out[84]
  PIN la_data_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9308 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.546 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1237.030000 0.000000 1237.170000 0.490000 ;
    END
  END la_data_out[83]
  PIN la_data_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9126 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.455 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1233.130000 0.000000 1233.270000 0.490000 ;
    END
  END la_data_out[82]
  PIN la_data_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9336 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.56 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1229.330000 0.000000 1229.470000 0.490000 ;
    END
  END la_data_out[81]
  PIN la_data_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1225.430000 0.000000 1225.570000 0.490000 ;
    END
  END la_data_out[80]
  PIN la_data_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8818 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.301 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1221.530000 0.000000 1221.670000 0.490000 ;
    END
  END la_data_out[79]
  PIN la_data_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9196 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.49 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1217.630000 0.000000 1217.770000 0.490000 ;
    END
  END la_data_out[78]
  PIN la_data_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1213.730000 0.000000 1213.870000 0.490000 ;
    END
  END la_data_out[77]
  PIN la_data_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1209.830000 0.000000 1209.970000 0.490000 ;
    END
  END la_data_out[76]
  PIN la_data_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.921 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.497 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1205.930000 0.000000 1206.070000 0.490000 ;
    END
  END la_data_out[75]
  PIN la_data_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9252 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.518 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1202.030000 0.000000 1202.170000 0.490000 ;
    END
  END la_data_out[74]
  PIN la_data_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1198.130000 0.000000 1198.270000 0.490000 ;
    END
  END la_data_out[73]
  PIN la_data_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.005 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.917 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1194.130000 0.000000 1194.270000 0.490000 ;
    END
  END la_data_out[72]
  PIN la_data_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9336 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.56 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1190.230000 0.000000 1190.370000 0.490000 ;
    END
  END la_data_out[71]
  PIN la_data_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1186.330000 0.000000 1186.470000 0.490000 ;
    END
  END la_data_out[70]
  PIN la_data_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9308 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.546 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1182.430000 0.000000 1182.570000 0.490000 ;
    END
  END la_data_out[69]
  PIN la_data_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.893 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.357 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1178.530000 0.000000 1178.670000 0.490000 ;
    END
  END la_data_out[68]
  PIN la_data_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.928 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.532 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1174.630000 0.000000 1174.770000 0.490000 ;
    END
  END la_data_out[67]
  PIN la_data_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9196 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.49 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1170.730000 0.000000 1170.870000 0.490000 ;
    END
  END la_data_out[66]
  PIN la_data_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8874 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.329 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1166.830000 0.000000 1166.970000 0.490000 ;
    END
  END la_data_out[65]
  PIN la_data_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1162.930000 0.000000 1163.070000 0.490000 ;
    END
  END la_data_out[64]
  PIN la_data_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9196 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.49 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1159.030000 0.000000 1159.170000 0.490000 ;
    END
  END la_data_out[63]
  PIN la_data_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.928 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.532 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1155.130000 0.000000 1155.270000 0.490000 ;
    END
  END la_data_out[62]
  PIN la_data_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.907 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.427 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1151.330000 0.000000 1151.470000 0.490000 ;
    END
  END la_data_out[61]
  PIN la_data_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1147.430000 0.000000 1147.570000 0.490000 ;
    END
  END la_data_out[60]
  PIN la_data_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1143.430000 0.000000 1143.570000 0.490000 ;
    END
  END la_data_out[59]
  PIN la_data_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9336 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.56 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1139.530000 0.000000 1139.670000 0.490000 ;
    END
  END la_data_out[58]
  PIN la_data_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1135.630000 0.000000 1135.770000 0.490000 ;
    END
  END la_data_out[57]
  PIN la_data_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9364 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.574 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1131.730000 0.000000 1131.870000 0.490000 ;
    END
  END la_data_out[56]
  PIN la_data_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1127.830000 0.000000 1127.970000 0.490000 ;
    END
  END la_data_out[55]
  PIN la_data_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8734 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.259 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1123.930000 0.000000 1124.070000 0.490000 ;
    END
  END la_data_out[54]
  PIN la_data_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1120.030000 0.000000 1120.170000 0.490000 ;
    END
  END la_data_out[53]
  PIN la_data_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.425 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.017 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1116.030000 0.000000 1116.170000 0.490000 ;
    END
  END la_data_out[52]
  PIN la_data_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9154 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.469 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1112.130000 0.000000 1112.270000 0.490000 ;
    END
  END la_data_out[51]
  PIN la_data_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1108.330000 0.000000 1108.470000 0.490000 ;
    END
  END la_data_out[50]
  PIN la_data_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1104.430000 0.000000 1104.570000 0.490000 ;
    END
  END la_data_out[49]
  PIN la_data_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1100.530000 0.000000 1100.670000 0.490000 ;
    END
  END la_data_out[48]
  PIN la_data_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8958 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.371 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1096.630000 0.000000 1096.770000 0.490000 ;
    END
  END la_data_out[47]
  PIN la_data_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9308 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.546 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1092.730000 0.000000 1092.870000 0.490000 ;
    END
  END la_data_out[46]
  PIN la_data_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1088.730000 0.000000 1088.870000 0.490000 ;
    END
  END la_data_out[45]
  PIN la_data_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9392 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.588 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1084.830000 0.000000 1084.970000 0.490000 ;
    END
  END la_data_out[44]
  PIN la_data_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1081.030000 0.000000 1081.170000 0.490000 ;
    END
  END la_data_out[43]
  PIN la_data_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9252 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.518 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1077.130000 0.000000 1077.270000 0.490000 ;
    END
  END la_data_out[42]
  PIN la_data_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9252 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.518 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1073.230000 0.000000 1073.370000 0.490000 ;
    END
  END la_data_out[41]
  PIN la_data_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8902 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1069.330000 0.000000 1069.470000 0.490000 ;
    END
  END la_data_out[40]
  PIN la_data_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1065.330000 0.000000 1065.470000 0.490000 ;
    END
  END la_data_out[39]
  PIN la_data_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1061.430000 0.000000 1061.570000 0.490000 ;
    END
  END la_data_out[38]
  PIN la_data_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1057.530000 0.000000 1057.670000 0.490000 ;
    END
  END la_data_out[37]
  PIN la_data_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9308 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.546 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1053.630000 0.000000 1053.770000 0.490000 ;
    END
  END la_data_out[36]
  PIN la_data_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1049.730000 0.000000 1049.870000 0.490000 ;
    END
  END la_data_out[35]
  PIN la_data_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1045.930000 0.000000 1046.070000 0.490000 ;
    END
  END la_data_out[34]
  PIN la_data_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9364 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.574 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1042.030000 0.000000 1042.170000 0.490000 ;
    END
  END la_data_out[33]
  PIN la_data_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1038.030000 0.000000 1038.170000 0.490000 ;
    END
  END la_data_out[32]
  PIN la_data_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9252 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.518 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1034.130000 0.000000 1034.270000 0.490000 ;
    END
  END la_data_out[31]
  PIN la_data_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9196 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.49 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1030.230000 0.000000 1030.370000 0.490000 ;
    END
  END la_data_out[30]
  PIN la_data_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.928 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.532 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1026.330000 0.000000 1026.470000 0.490000 ;
    END
  END la_data_out[29]
  PIN la_data_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9196 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.49 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1022.430000 0.000000 1022.570000 0.490000 ;
    END
  END la_data_out[28]
  PIN la_data_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9308 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.546 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1018.530000 0.000000 1018.670000 0.490000 ;
    END
  END la_data_out[27]
  PIN la_data_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1014.630000 0.000000 1014.770000 0.490000 ;
    END
  END la_data_out[26]
  PIN la_data_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9336 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.56 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1010.730000 0.000000 1010.870000 0.490000 ;
    END
  END la_data_out[25]
  PIN la_data_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1006.830000 0.000000 1006.970000 0.490000 ;
    END
  END la_data_out[24]
  PIN la_data_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1002.930000 0.000000 1003.070000 0.490000 ;
    END
  END la_data_out[23]
  PIN la_data_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9966 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.875 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 999.030000 0.000000 999.170000 0.490000 ;
    END
  END la_data_out[22]
  PIN la_data_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 995.130000 0.000000 995.270000 0.490000 ;
    END
  END la_data_out[21]
  PIN la_data_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.413 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 991.230000 0.000000 991.370000 0.490000 ;
    END
  END la_data_out[20]
  PIN la_data_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.935 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.567 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 987.330000 0.000000 987.470000 0.490000 ;
    END
  END la_data_out[19]
  PIN la_data_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9014 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.399 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 983.430000 0.000000 983.570000 0.490000 ;
    END
  END la_data_out[18]
  PIN la_data_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9322 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.553 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 979.530000 0.000000 979.670000 0.490000 ;
    END
  END la_data_out[17]
  PIN la_data_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9098 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.441 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 975.630000 0.000000 975.770000 0.490000 ;
    END
  END la_data_out[16]
  PIN la_data_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.879 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.287 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 971.730000 0.000000 971.870000 0.490000 ;
    END
  END la_data_out[15]
  PIN la_data_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9126 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.455 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 967.830000 0.000000 967.970000 0.490000 ;
    END
  END la_data_out[14]
  PIN la_data_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9266 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.525 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 963.930000 0.000000 964.070000 0.490000 ;
    END
  END la_data_out[13]
  PIN la_data_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9014 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.399 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 959.930000 0.000000 960.070000 0.490000 ;
    END
  END la_data_out[12]
  PIN la_data_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.935 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.567 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 956.030000 0.000000 956.170000 0.490000 ;
    END
  END la_data_out[11]
  PIN la_data_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.413 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 952.130000 0.000000 952.270000 0.490000 ;
    END
  END la_data_out[10]
  PIN la_data_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.935 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.567 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 948.230000 0.000000 948.370000 0.490000 ;
    END
  END la_data_out[9]
  PIN la_data_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9014 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.399 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 944.330000 0.000000 944.470000 0.490000 ;
    END
  END la_data_out[8]
  PIN la_data_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9322 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.553 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 940.430000 0.000000 940.570000 0.490000 ;
    END
  END la_data_out[7]
  PIN la_data_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9238 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.511 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 936.630000 0.000000 936.770000 0.490000 ;
    END
  END la_data_out[6]
  PIN la_data_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 932.630000 0.000000 932.770000 0.490000 ;
    END
  END la_data_out[5]
  PIN la_data_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9126 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.455 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 928.730000 0.000000 928.870000 0.490000 ;
    END
  END la_data_out[4]
  PIN la_data_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9126 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.455 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 924.930000 0.000000 925.070000 0.490000 ;
    END
  END la_data_out[3]
  PIN la_data_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 921.030000 0.000000 921.170000 0.490000 ;
    END
  END la_data_out[2]
  PIN la_data_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9098 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.441 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 917.130000 0.000000 917.270000 0.490000 ;
    END
  END la_data_out[1]
  PIN la_data_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8762 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.273 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 913.230000 0.000000 913.370000 0.490000 ;
    END
  END la_data_out[0]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1908.530000 0.000000 1908.670000 0.490000 ;
    END
  END la_oenb[127]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1904.630000 0.000000 1904.770000 0.490000 ;
    END
  END la_oenb[126]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1900.730000 0.000000 1900.870000 0.490000 ;
    END
  END la_oenb[125]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1896.730000 0.000000 1896.870000 0.490000 ;
    END
  END la_oenb[124]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1892.830000 0.000000 1892.970000 0.490000 ;
    END
  END la_oenb[123]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1888.930000 0.000000 1889.070000 0.490000 ;
    END
  END la_oenb[122]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1885.030000 0.000000 1885.170000 0.490000 ;
    END
  END la_oenb[121]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1881.130000 0.000000 1881.270000 0.490000 ;
    END
  END la_oenb[120]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1877.230000 0.000000 1877.370000 0.490000 ;
    END
  END la_oenb[119]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1873.330000 0.000000 1873.470000 0.490000 ;
    END
  END la_oenb[118]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1869.430000 0.000000 1869.570000 0.490000 ;
    END
  END la_oenb[117]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1865.530000 0.000000 1865.670000 0.490000 ;
    END
  END la_oenb[116]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1861.630000 0.000000 1861.770000 0.490000 ;
    END
  END la_oenb[115]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1857.730000 0.000000 1857.870000 0.490000 ;
    END
  END la_oenb[114]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1853.830000 0.000000 1853.970000 0.490000 ;
    END
  END la_oenb[113]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1849.930000 0.000000 1850.070000 0.490000 ;
    END
  END la_oenb[112]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1846.030000 0.000000 1846.170000 0.490000 ;
    END
  END la_oenb[111]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1842.130000 0.000000 1842.270000 0.490000 ;
    END
  END la_oenb[110]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1838.230000 0.000000 1838.370000 0.490000 ;
    END
  END la_oenb[109]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1834.330000 0.000000 1834.470000 0.490000 ;
    END
  END la_oenb[108]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1830.430000 0.000000 1830.570000 0.490000 ;
    END
  END la_oenb[107]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1826.530000 0.000000 1826.670000 0.490000 ;
    END
  END la_oenb[106]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1822.630000 0.000000 1822.770000 0.490000 ;
    END
  END la_oenb[105]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1818.630000 0.000000 1818.770000 0.490000 ;
    END
  END la_oenb[104]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1814.730000 0.000000 1814.870000 0.490000 ;
    END
  END la_oenb[103]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1810.830000 0.000000 1810.970000 0.490000 ;
    END
  END la_oenb[102]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1806.930000 0.000000 1807.070000 0.490000 ;
    END
  END la_oenb[101]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1803.030000 0.000000 1803.170000 0.490000 ;
    END
  END la_oenb[100]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1799.230000 0.000000 1799.370000 0.490000 ;
    END
  END la_oenb[99]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1795.330000 0.000000 1795.470000 0.490000 ;
    END
  END la_oenb[98]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1791.330000 0.000000 1791.470000 0.490000 ;
    END
  END la_oenb[97]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1787.530000 0.000000 1787.670000 0.490000 ;
    END
  END la_oenb[96]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1783.630000 0.000000 1783.770000 0.490000 ;
    END
  END la_oenb[95]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1779.730000 0.000000 1779.870000 0.490000 ;
    END
  END la_oenb[94]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1775.830000 0.000000 1775.970000 0.490000 ;
    END
  END la_oenb[93]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1771.930000 0.000000 1772.070000 0.490000 ;
    END
  END la_oenb[92]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1767.930000 0.000000 1768.070000 0.490000 ;
    END
  END la_oenb[91]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1764.030000 0.000000 1764.170000 0.490000 ;
    END
  END la_oenb[90]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1760.130000 0.000000 1760.270000 0.490000 ;
    END
  END la_oenb[89]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1756.230000 0.000000 1756.370000 0.490000 ;
    END
  END la_oenb[88]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1752.330000 0.000000 1752.470000 0.490000 ;
    END
  END la_oenb[87]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1748.430000 0.000000 1748.570000 0.490000 ;
    END
  END la_oenb[86]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1744.530000 0.000000 1744.670000 0.490000 ;
    END
  END la_oenb[85]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1740.530000 0.000000 1740.670000 0.490000 ;
    END
  END la_oenb[84]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1736.630000 0.000000 1736.770000 0.490000 ;
    END
  END la_oenb[83]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1732.730000 0.000000 1732.870000 0.490000 ;
    END
  END la_oenb[82]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1728.930000 0.000000 1729.070000 0.490000 ;
    END
  END la_oenb[81]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1725.030000 0.000000 1725.170000 0.490000 ;
    END
  END la_oenb[80]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1721.230000 0.000000 1721.370000 0.490000 ;
    END
  END la_oenb[79]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1717.330000 0.000000 1717.470000 0.490000 ;
    END
  END la_oenb[78]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1713.330000 0.000000 1713.470000 0.490000 ;
    END
  END la_oenb[77]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1709.430000 0.000000 1709.570000 0.490000 ;
    END
  END la_oenb[76]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1705.530000 0.000000 1705.670000 0.490000 ;
    END
  END la_oenb[75]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1701.630000 0.000000 1701.770000 0.490000 ;
    END
  END la_oenb[74]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1697.730000 0.000000 1697.870000 0.490000 ;
    END
  END la_oenb[73]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1693.830000 0.000000 1693.970000 0.490000 ;
    END
  END la_oenb[72]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1689.830000 0.000000 1689.970000 0.490000 ;
    END
  END la_oenb[71]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1685.930000 0.000000 1686.070000 0.490000 ;
    END
  END la_oenb[70]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1682.030000 0.000000 1682.170000 0.490000 ;
    END
  END la_oenb[69]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1678.130000 0.000000 1678.270000 0.490000 ;
    END
  END la_oenb[68]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1674.230000 0.000000 1674.370000 0.490000 ;
    END
  END la_oenb[67]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1670.330000 0.000000 1670.470000 0.490000 ;
    END
  END la_oenb[66]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1666.430000 0.000000 1666.570000 0.490000 ;
    END
  END la_oenb[65]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1662.530000 0.000000 1662.670000 0.490000 ;
    END
  END la_oenb[64]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1658.630000 0.000000 1658.770000 0.490000 ;
    END
  END la_oenb[63]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1654.830000 0.000000 1654.970000 0.490000 ;
    END
  END la_oenb[62]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1650.930000 0.000000 1651.070000 0.490000 ;
    END
  END la_oenb[61]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1647.030000 0.000000 1647.170000 0.490000 ;
    END
  END la_oenb[60]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1643.130000 0.000000 1643.270000 0.490000 ;
    END
  END la_oenb[59]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1639.230000 0.000000 1639.370000 0.490000 ;
    END
  END la_oenb[58]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1635.230000 0.000000 1635.370000 0.490000 ;
    END
  END la_oenb[57]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1631.330000 0.000000 1631.470000 0.490000 ;
    END
  END la_oenb[56]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1627.430000 0.000000 1627.570000 0.490000 ;
    END
  END la_oenb[55]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1623.530000 0.000000 1623.670000 0.490000 ;
    END
  END la_oenb[54]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1619.630000 0.000000 1619.770000 0.490000 ;
    END
  END la_oenb[53]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1615.730000 0.000000 1615.870000 0.490000 ;
    END
  END la_oenb[52]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1611.730000 0.000000 1611.870000 0.490000 ;
    END
  END la_oenb[51]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1607.830000 0.000000 1607.970000 0.490000 ;
    END
  END la_oenb[50]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1603.930000 0.000000 1604.070000 0.490000 ;
    END
  END la_oenb[49]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1600.130000 0.000000 1600.270000 0.490000 ;
    END
  END la_oenb[48]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1596.230000 0.000000 1596.370000 0.490000 ;
    END
  END la_oenb[47]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1592.330000 0.000000 1592.470000 0.490000 ;
    END
  END la_oenb[46]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1588.430000 0.000000 1588.570000 0.490000 ;
    END
  END la_oenb[45]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1584.530000 0.000000 1584.670000 0.490000 ;
    END
  END la_oenb[44]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1580.630000 0.000000 1580.770000 0.490000 ;
    END
  END la_oenb[43]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1576.730000 0.000000 1576.870000 0.490000 ;
    END
  END la_oenb[42]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1572.830000 0.000000 1572.970000 0.490000 ;
    END
  END la_oenb[41]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1568.930000 0.000000 1569.070000 0.490000 ;
    END
  END la_oenb[40]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1565.030000 0.000000 1565.170000 0.490000 ;
    END
  END la_oenb[39]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1561.130000 0.000000 1561.270000 0.490000 ;
    END
  END la_oenb[38]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1557.130000 0.000000 1557.270000 0.490000 ;
    END
  END la_oenb[37]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1553.230000 0.000000 1553.370000 0.490000 ;
    END
  END la_oenb[36]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1549.330000 0.000000 1549.470000 0.490000 ;
    END
  END la_oenb[35]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1545.430000 0.000000 1545.570000 0.490000 ;
    END
  END la_oenb[34]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1541.530000 0.000000 1541.670000 0.490000 ;
    END
  END la_oenb[33]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1537.730000 0.000000 1537.870000 0.490000 ;
    END
  END la_oenb[32]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1533.730000 0.000000 1533.870000 0.490000 ;
    END
  END la_oenb[31]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1529.830000 0.000000 1529.970000 0.490000 ;
    END
  END la_oenb[30]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1525.930000 0.000000 1526.070000 0.490000 ;
    END
  END la_oenb[29]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1522.030000 0.000000 1522.170000 0.490000 ;
    END
  END la_oenb[28]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1518.130000 0.000000 1518.270000 0.490000 ;
    END
  END la_oenb[27]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1514.230000 0.000000 1514.370000 0.490000 ;
    END
  END la_oenb[26]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1510.430000 0.000000 1510.570000 0.490000 ;
    END
  END la_oenb[25]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1506.430000 0.000000 1506.570000 0.490000 ;
    END
  END la_oenb[24]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1502.530000 0.000000 1502.670000 0.490000 ;
    END
  END la_oenb[23]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1498.630000 0.000000 1498.770000 0.490000 ;
    END
  END la_oenb[22]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1494.730000 0.000000 1494.870000 0.490000 ;
    END
  END la_oenb[21]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1490.830000 0.000000 1490.970000 0.490000 ;
    END
  END la_oenb[20]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1486.930000 0.000000 1487.070000 0.490000 ;
    END
  END la_oenb[19]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1483.030000 0.000000 1483.170000 0.490000 ;
    END
  END la_oenb[18]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1479.130000 0.000000 1479.270000 0.490000 ;
    END
  END la_oenb[17]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1475.230000 0.000000 1475.370000 0.490000 ;
    END
  END la_oenb[16]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1471.330000 0.000000 1471.470000 0.490000 ;
    END
  END la_oenb[15]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1467.430000 0.000000 1467.570000 0.490000 ;
    END
  END la_oenb[14]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1463.530000 0.000000 1463.670000 0.490000 ;
    END
  END la_oenb[13]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1459.630000 0.000000 1459.770000 0.490000 ;
    END
  END la_oenb[12]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1455.630000 0.000000 1455.770000 0.490000 ;
    END
  END la_oenb[11]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1451.730000 0.000000 1451.870000 0.490000 ;
    END
  END la_oenb[10]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1447.830000 0.000000 1447.970000 0.490000 ;
    END
  END la_oenb[9]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1443.930000 0.000000 1444.070000 0.490000 ;
    END
  END la_oenb[8]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1440.130000 0.000000 1440.270000 0.490000 ;
    END
  END la_oenb[7]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1436.230000 0.000000 1436.370000 0.490000 ;
    END
  END la_oenb[6]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1432.330000 0.000000 1432.470000 0.490000 ;
    END
  END la_oenb[5]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1428.330000 0.000000 1428.470000 0.490000 ;
    END
  END la_oenb[4]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1424.430000 0.000000 1424.570000 0.490000 ;
    END
  END la_oenb[3]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1420.530000 0.000000 1420.670000 0.490000 ;
    END
  END la_oenb[2]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1416.730000 0.000000 1416.870000 0.490000 ;
    END
  END la_oenb[1]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1412.830000 0.000000 1412.970000 0.490000 ;
    END
  END la_oenb[0]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 94.890000 0.800000 95.190000 ;
    END
  END io_in[37]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8788 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.152 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.9618 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 21.6 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 43.1336 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 211.717 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 237.835000 0.800000 238.135000 ;
    END
  END io_in[36]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 93.0316 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 496.16 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.318 LAYER met4  ;
    ANTENNAMAXAREACAR 23.989 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 122.601 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.413208 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 380.780000 0.800000 381.080000 ;
    END
  END io_in[35]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 571.530000 0.800000 571.830000 ;
    END
  END io_in[34]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.8919 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 53.2 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.1448 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.576 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 31.5399 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 167.918 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 761.995000 0.800000 762.295000 ;
    END
  END io_in[33]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 177.903 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 949.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 76.6032 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 410.432 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 150.942 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 791.152 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.208175 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 952.650000 0.800000 952.950000 ;
    END
  END io_in[32]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2843 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.3758 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 23.808 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 22.0808 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 110.399 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.460202 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1143.500000 0.800000 1143.800000 ;
    END
  END io_in[31]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2909 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.328 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.3758 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 23.808 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met4  ;
    ANTENNAMAXAREACAR 11.5846 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 56.284 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.381719 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1333.865000 0.800000 1334.165000 ;
    END
  END io_in[30]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4803 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.36 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.1448 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.576 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 32.312 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 168.941 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1524.520000 0.800000 1524.820000 ;
    END
  END io_in[29]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.6082 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3534 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.88 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8047 LAYER met3  ;
    ANTENNAMAXAREACAR 82.1173 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 389.309 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.169358 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1715.180000 0.800000 1715.480000 ;
    END
  END io_in[28]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1308 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.496 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.1448 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.576 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 38.6763 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 201.964 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1905.835000 0.800000 1906.135000 ;
    END
  END io_in[27]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 110.238 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 588.4 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 62.1865 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 316.843 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2096.490000 0.800000 2096.790000 ;
    END
  END io_in[26]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.1735 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.6149 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.608 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.3325 LAYER met3  ;
    ANTENNAMAXAREACAR 83.9677 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 402.878 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.135391 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2287.145000 0.800000 2287.445000 ;
    END
  END io_in[25]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 107.603 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 574.344 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 19.1884 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 104.377 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2477.705000 0.800000 2478.005000 ;
    END
  END io_in[24]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.730000 2594.730000 109.870000 2595.220000 ;
    END
  END io_in[23]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.630000 2594.730000 329.770000 2595.220000 ;
    END
  END io_in[22]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.530000 2594.730000 549.670000 2595.220000 ;
    END
  END io_in[21]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.430000 2594.730000 769.570000 2595.220000 ;
    END
  END io_in[20]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 989.430000 2594.730000 989.570000 2595.220000 ;
    END
  END io_in[19]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1209.330000 2594.730000 1209.470000 2595.220000 ;
    END
  END io_in[18]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1429.230000 2594.730000 1429.370000 2595.220000 ;
    END
  END io_in[17]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1649.130000 2594.730000 1649.270000 2595.220000 ;
    END
  END io_in[16]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1869.130000 2594.730000 1869.270000 2595.220000 ;
    END
  END io_in[15]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 2428.265000 1926.480000 2428.565000 ;
    END
  END io_in[14]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 2233.865000 1926.480000 2234.165000 ;
    END
  END io_in[13]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 2039.660000 1926.480000 2039.960000 ;
    END
  END io_in[12]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 1845.355000 1926.480000 1845.655000 ;
    END
  END io_in[11]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 1651.050000 1926.480000 1651.350000 ;
    END
  END io_in[10]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 1456.840000 1926.480000 1457.140000 ;
    END
  END io_in[9]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 77.0688 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 412.888 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.139 LAYER met3  ;
    ANTENNAMAXAREACAR 62.7292 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 323.781 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.445596 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.1708 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 44.048 LAYER met4  ;
    ANTENNAGATEAREA 2.3355 LAYER met4  ;
    ANTENNAMAXAREACAR 66.2277 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 342.641 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 1262.440000 1926.480000 1262.740000 ;
    END
  END io_in[8]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 1068.140000 1926.480000 1068.440000 ;
    END
  END io_in[7]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 873.930000 1926.480000 874.230000 ;
    END
  END io_in[6]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0546 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.616 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 45.3918 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 242.56 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 101.204 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 517.655 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.208175 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 728.300000 1926.480000 728.600000 ;
    END
  END io_in[5]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 582.475000 1926.480000 582.775000 ;
    END
  END io_in[4]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 436.745000 1926.480000 437.045000 ;
    END
  END io_in[3]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 291.115000 1926.480000 291.415000 ;
    END
  END io_in[2]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 145.385000 1926.480000 145.685000 ;
    END
  END io_in[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 1.865000 1926.480000 2.165000 ;
    END
  END io_in[0]
  PIN io_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 37.9363 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 202.792 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.7918 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 31.36 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 48.8588 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 257.415 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 47.180000 0.800000 47.480000 ;
    END
  END io_out[37]
  PIN io_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3354 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.784 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 190.120000 0.800000 190.420000 ;
    END
  END io_out[36]
  PIN io_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0964 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.176 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 333.160000 0.800000 333.460000 ;
    END
  END io_out[35]
  PIN io_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 131.997 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 704.448 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 61.2888 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 327.344 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 523.820000 0.800000 524.120000 ;
    END
  END io_out[34]
  PIN io_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.872 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 714.475000 0.800000 714.775000 ;
    END
  END io_out[33]
  PIN io_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.872 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 904.940000 0.800000 905.240000 ;
    END
  END io_out[32]
  PIN io_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.872 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1095.785000 0.800000 1096.085000 ;
    END
  END io_out[31]
  PIN io_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.872 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1286.250000 0.800000 1286.550000 ;
    END
  END io_out[30]
  PIN io_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.872 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1476.810000 0.800000 1477.110000 ;
    END
  END io_out[29]
  PIN io_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9264 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.936 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1667.660000 0.800000 1667.960000 ;
    END
  END io_out[28]
  PIN io_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3174 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.688 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1858.220000 0.800000 1858.520000 ;
    END
  END io_out[27]
  PIN io_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.0994 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.192 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2048.680000 0.800000 2048.980000 ;
    END
  END io_out[26]
  PIN io_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2499 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2239.435000 0.800000 2239.735000 ;
    END
  END io_out[25]
  PIN io_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1989 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.056 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2430.185000 0.800000 2430.485000 ;
    END
  END io_out[24]
  PIN io_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.11 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.442 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 54.830000 2594.730000 54.970000 2595.220000 ;
    END
  END io_out[23]
  PIN io_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.11 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.442 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 274.630000 2594.730000 274.770000 2595.220000 ;
    END
  END io_out[22]
  PIN io_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.11 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.442 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 494.530000 2594.730000 494.670000 2595.220000 ;
    END
  END io_out[21]
  PIN io_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.11 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.442 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 714.430000 2594.730000 714.570000 2595.220000 ;
    END
  END io_out[20]
  PIN io_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.268 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.114 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 934.530000 2594.730000 934.670000 2595.220000 ;
    END
  END io_out[19]
  PIN io_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2582 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.065 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1154.430000 2594.730000 1154.570000 2595.220000 ;
    END
  END io_out[18]
  PIN io_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.1808 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.7982 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.765 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1374.330000 2594.730000 1374.470000 2595.220000 ;
    END
  END io_out[17]
  PIN io_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.1808 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.38 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.792 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1594.230000 2594.730000 1594.370000 2595.220000 ;
    END
  END io_out[16]
  PIN io_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 74.4791 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 372.117 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.3768 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 98.48 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1814.230000 2594.730000 1814.370000 2595.220000 ;
    END
  END io_out[15]
  PIN io_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4404 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.344 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 2476.840000 1926.480000 2477.140000 ;
    END
  END io_out[14]
  PIN io_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7334 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 2282.440000 1926.480000 2282.740000 ;
    END
  END io_out[13]
  PIN io_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 2088.140000 1926.480000 2088.440000 ;
    END
  END io_out[12]
  PIN io_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3444 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.832 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 1894.120000 1926.480000 1894.420000 ;
    END
  END io_out[11]
  PIN io_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5784 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.08 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 1699.720000 1926.480000 1700.020000 ;
    END
  END io_out[10]
  PIN io_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.1874 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 38.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 1505.320000 1926.480000 1505.620000 ;
    END
  END io_out[9]
  PIN io_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3764 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.336 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 1311.020000 1926.480000 1311.320000 ;
    END
  END io_out[8]
  PIN io_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3849 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.048 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 1116.715000 1926.480000 1117.015000 ;
    END
  END io_out[7]
  PIN io_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.472 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 922.410000 1926.480000 922.710000 ;
    END
  END io_out[6]
  PIN io_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4404 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.344 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 776.680000 1926.480000 776.980000 ;
    END
  END io_out[5]
  PIN io_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5062 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.832 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 631.050000 1926.480000 631.350000 ;
    END
  END io_out[4]
  PIN io_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6069 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.232 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 485.225000 1926.480000 485.525000 ;
    END
  END io_out[3]
  PIN io_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3596 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.616 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 11.6478 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 62.592 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 339.500000 1926.480000 339.800000 ;
    END
  END io_out[2]
  PIN io_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6489 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.456 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 193.865000 1926.480000 194.165000 ;
    END
  END io_out[1]
  PIN io_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.872 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 47.945000 1926.480000 48.245000 ;
    END
  END io_out[0]
  PIN io_oeb[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3624 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.928 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 0.620000 0.800000 0.920000 ;
    END
  END io_oeb[37]
  PIN io_oeb[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4029 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.144 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 142.505000 0.800000 142.805000 ;
    END
  END io_oeb[36]
  PIN io_oeb[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5244 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.792 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 285.450000 0.800000 285.750000 ;
    END
  END io_oeb[35]
  PIN io_oeb[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.872 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 476.010000 0.800000 476.310000 ;
    END
  END io_oeb[34]
  PIN io_oeb[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.872 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 666.860000 0.800000 667.160000 ;
    END
  END io_oeb[33]
  PIN io_oeb[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.872 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 857.320000 0.800000 857.620000 ;
    END
  END io_oeb[32]
  PIN io_oeb[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5154 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.744 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1047.980000 0.800000 1048.280000 ;
    END
  END io_oeb[31]
  PIN io_oeb[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7664 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.416 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1238.730000 0.800000 1239.030000 ;
    END
  END io_oeb[30]
  PIN io_oeb[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.0009 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1429.195000 0.800000 1429.495000 ;
    END
  END io_oeb[29]
  PIN io_oeb[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.8719 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.312 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1619.945000 0.800000 1620.245000 ;
    END
  END io_oeb[28]
  PIN io_oeb[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2199 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.168 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1810.505000 0.800000 1810.805000 ;
    END
  END io_oeb[27]
  PIN io_oeb[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3204 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.704 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2001.160000 0.800000 2001.460000 ;
    END
  END io_oeb[26]
  PIN io_oeb[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2394 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.272 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2191.820000 0.800000 2192.120000 ;
    END
  END io_oeb[25]
  PIN io_oeb[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8727 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2382.475000 0.800000 2382.775000 ;
    END
  END io_oeb[24]
  PIN io_oeb[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1107 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.4455 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 3.630000 2594.735000 3.770000 2595.220000 ;
    END
  END io_oeb[23]
  PIN io_oeb[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.11 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.442 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 219.730000 2594.730000 219.870000 2595.220000 ;
    END
  END io_oeb[22]
  PIN io_oeb[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.11 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.442 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 439.630000 2594.730000 439.770000 2595.220000 ;
    END
  END io_oeb[21]
  PIN io_oeb[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.11 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.442 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 659.530000 2594.730000 659.670000 2595.220000 ;
    END
  END io_oeb[20]
  PIN io_oeb[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6348 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.066 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 879.530000 2594.730000 879.670000 2595.220000 ;
    END
  END io_oeb[19]
  PIN io_oeb[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3212 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.498 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1099.430000 2594.730000 1099.570000 2595.220000 ;
    END
  END io_oeb[18]
  PIN io_oeb[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 73.9232 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 369.39 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1319.330000 2594.730000 1319.470000 2595.220000 ;
    END
  END io_oeb[17]
  PIN io_oeb[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.1808 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.107 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.427 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1539.230000 2594.730000 1539.370000 2595.220000 ;
    END
  END io_oeb[16]
  PIN io_oeb[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6207 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.8035 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.2968 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 60.72 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1759.230000 2594.730000 1759.370000 2595.220000 ;
    END
  END io_oeb[15]
  PIN io_oeb[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3444 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.832 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 2523.400000 1926.480000 2523.700000 ;
    END
  END io_oeb[14]
  PIN io_oeb[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3269 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.072 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 2331.115000 1926.480000 2331.415000 ;
    END
  END io_oeb[13]
  PIN io_oeb[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4314 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.296 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 2136.810000 1926.480000 2137.110000 ;
    END
  END io_oeb[12]
  PIN io_oeb[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.3699 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.968 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 1942.505000 1926.480000 1942.805000 ;
    END
  END io_oeb[11]
  PIN io_oeb[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3774 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.008 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 1748.200000 1926.480000 1748.500000 ;
    END
  END io_oeb[10]
  PIN io_oeb[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2679 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.424 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 1553.995000 1926.480000 1554.295000 ;
    END
  END io_oeb[9]
  PIN io_oeb[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7036 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.744 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 80.6466 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 431.056 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 1359.690000 1926.480000 1359.990000 ;
    END
  END io_oeb[8]
  PIN io_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2979 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 1165.385000 1926.480000 1165.685000 ;
    END
  END io_oeb[7]
  PIN io_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2229 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 970.985000 1926.480000 971.285000 ;
    END
  END io_oeb[6]
  PIN io_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4139 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.536 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 825.355000 1926.480000 825.655000 ;
    END
  END io_oeb[5]
  PIN io_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5259 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.8 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 679.625000 1926.480000 679.925000 ;
    END
  END io_oeb[4]
  PIN io_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.096 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 533.900000 1926.480000 534.200000 ;
    END
  END io_oeb[3]
  PIN io_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0149 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.408 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 388.075000 1926.480000 388.375000 ;
    END
  END io_oeb[2]
  PIN io_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.36235 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.624 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 22.8108 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 122.128 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 242.345000 1926.480000 242.645000 ;
    END
  END io_oeb[1]
  PIN io_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6121 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.256 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.8898 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 37.216 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 96.715000 1926.480000 97.015000 ;
    END
  END io_oeb[0]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 428.490000 0.800000 428.790000 ;
    END
  END analog_io[28]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 619.145000 0.800000 619.445000 ;
    END
  END analog_io[27]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 809.610000 0.800000 809.910000 ;
    END
  END analog_io[26]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1000.265000 0.800000 1000.565000 ;
    END
  END analog_io[25]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1191.020000 0.800000 1191.320000 ;
    END
  END analog_io[24]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1381.580000 0.800000 1381.880000 ;
    END
  END analog_io[23]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1572.330000 0.800000 1572.630000 ;
    END
  END analog_io[22]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1762.890000 0.800000 1763.190000 ;
    END
  END analog_io[21]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1953.450000 0.800000 1953.750000 ;
    END
  END analog_io[20]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2144.105000 0.800000 2144.405000 ;
    END
  END analog_io[19]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2334.665000 0.800000 2334.965000 ;
    END
  END analog_io[18]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2522.825000 0.800000 2523.125000 ;
    END
  END analog_io[17]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.730000 2594.730000 164.870000 2595.220000 ;
    END
  END analog_io[16]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.630000 2594.730000 384.770000 2595.220000 ;
    END
  END analog_io[15]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.530000 2594.730000 604.670000 2595.220000 ;
    END
  END analog_io[14]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.530000 2594.730000 824.670000 2595.220000 ;
    END
  END analog_io[13]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1044.430000 2594.730000 1044.570000 2595.220000 ;
    END
  END analog_io[12]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1264.330000 2594.730000 1264.470000 2595.220000 ;
    END
  END analog_io[11]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1484.230000 2594.730000 1484.370000 2595.220000 ;
    END
  END analog_io[10]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1704.230000 2594.730000 1704.370000 2595.220000 ;
    END
  END analog_io[9]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1921.030000 2594.735000 1921.170000 2595.220000 ;
    END
  END analog_io[8]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 2379.785000 1926.480000 2380.085000 ;
    END
  END analog_io[7]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 2185.385000 1926.480000 2185.685000 ;
    END
  END analog_io[6]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 1991.080000 1926.480000 1991.380000 ;
    END
  END analog_io[5]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 1796.780000 1926.480000 1797.080000 ;
    END
  END analog_io[4]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 1602.380000 1926.480000 1602.680000 ;
    END
  END analog_io[3]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 1408.075000 1926.480000 1408.375000 ;
    END
  END analog_io[2]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 1214.060000 1926.480000 1214.360000 ;
    END
  END analog_io[1]
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1925.680000 1019.660000 1926.480000 1019.960000 ;
    END
  END analog_io[0]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1912.330000 0.000000 1912.470000 0.490000 ;
    END
  END user_clock2
  PIN user_irq[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9735 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.7595 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1922.730000 0.000000 1922.870000 0.485000 ;
    END
  END user_irq[2]
  PIN user_irq[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0874 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.211 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1920.130000 0.000000 1920.270000 0.490000 ;
    END
  END user_irq[1]
  PIN user_irq[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9672 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.728 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1916.230000 0.000000 1916.370000 0.490000 ;
    END
  END user_irq[0]
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 6.980000 7.260000 1919.500000 11.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.980000 2582.940000 1919.500000 2586.940000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1915.500000 7.260000 1919.500000 2586.940000 ;
    END
    PORT
      LAYER met4 ;
        RECT 6.980000 7.260000 10.980000 2586.940000 ;
    END

# P/G pin shape extracted from block 'tcam_32x28'
    PORT
      LAYER met4 ;
        RECT 824.905000 2125.920000 826.645000 2520.700000 ;
      LAYER met3 ;
        RECT 824.905000 2518.960000 1301.965000 2520.700000 ;
      LAYER met3 ;
        RECT 824.905000 2125.920000 1301.965000 2127.660000 ;
      LAYER met4 ;
        RECT 1300.225000 2125.920000 1301.965000 2520.700000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1387.045000 2126.015000 1388.785000 2520.795000 ;
      LAYER met3 ;
        RECT 1387.045000 2519.055000 1864.105000 2520.795000 ;
      LAYER met3 ;
        RECT 1387.045000 2126.015000 1864.105000 2127.755000 ;
      LAYER met4 ;
        RECT 1862.365000 2126.015000 1864.105000 2520.795000 ;
    END
    PORT
      LAYER met4 ;
        RECT 798.835000 2086.485000 800.835000 2556.325000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1888.375000 2086.485000 1890.375000 2556.325000 ;
    END
    PORT
      LAYER met3 ;
        RECT 798.835000 2554.325000 1890.375000 2556.325000 ;
    END
    PORT
      LAYER met3 ;
        RECT 798.835000 2086.485000 1890.375000 2088.485000 ;
    END
# end of P/G pin shape extracted from block 'tcam_32x28'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1897.460000 83.190000 1899.200000 477.970000 ;
      LAYER met3 ;
        RECT 1422.140000 83.190000 1899.200000 84.930000 ;
      LAYER met3 ;
        RECT 1422.140000 476.230000 1899.200000 477.970000 ;
      LAYER met4 ;
        RECT 1422.140000 83.190000 1423.880000 477.970000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1897.460000 592.890000 1899.200000 987.670000 ;
      LAYER met3 ;
        RECT 1422.140000 592.890000 1899.200000 594.630000 ;
      LAYER met3 ;
        RECT 1422.140000 985.930000 1899.200000 987.670000 ;
      LAYER met4 ;
        RECT 1422.140000 592.890000 1423.880000 987.670000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1897.460000 1102.590000 1899.200000 1497.370000 ;
      LAYER met3 ;
        RECT 1422.140000 1102.590000 1899.200000 1104.330000 ;
      LAYER met3 ;
        RECT 1422.140000 1495.630000 1899.200000 1497.370000 ;
      LAYER met4 ;
        RECT 1422.140000 1102.590000 1423.880000 1497.370000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1897.460000 1612.290000 1899.200000 2007.070000 ;
      LAYER met3 ;
        RECT 1422.140000 1612.290000 1899.200000 1614.030000 ;
      LAYER met3 ;
        RECT 1422.140000 2005.330000 1899.200000 2007.070000 ;
      LAYER met4 ;
        RECT 1422.140000 1612.290000 1423.880000 2007.070000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1264.680000 83.190000 1266.420000 477.970000 ;
      LAYER met3 ;
        RECT 789.360000 83.190000 1266.420000 84.930000 ;
      LAYER met3 ;
        RECT 789.360000 476.230000 1266.420000 477.970000 ;
      LAYER met4 ;
        RECT 789.360000 83.190000 791.100000 477.970000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1264.680000 592.890000 1266.420000 987.670000 ;
      LAYER met3 ;
        RECT 789.360000 592.890000 1266.420000 594.630000 ;
      LAYER met3 ;
        RECT 789.360000 985.930000 1266.420000 987.670000 ;
      LAYER met4 ;
        RECT 789.360000 592.890000 791.100000 987.670000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1264.680000 1102.590000 1266.420000 1497.370000 ;
      LAYER met3 ;
        RECT 789.360000 1102.590000 1266.420000 1104.330000 ;
      LAYER met3 ;
        RECT 789.360000 1495.630000 1266.420000 1497.370000 ;
      LAYER met4 ;
        RECT 789.360000 1102.590000 791.100000 1497.370000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1264.680000 1612.290000 1266.420000 2007.070000 ;
      LAYER met3 ;
        RECT 789.360000 1612.290000 1266.420000 1614.030000 ;
      LAYER met3 ;
        RECT 789.360000 2005.330000 1266.420000 2007.070000 ;
      LAYER met4 ;
        RECT 789.360000 1612.290000 791.100000 2007.070000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END vssd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 12.780000 2577.140000 1913.700000 2581.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.780000 13.060000 1913.700000 17.060000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1909.700000 13.060000 1913.700000 2581.140000 ;
    END
    PORT
      LAYER met4 ;
        RECT 12.780000 13.060000 16.780000 2581.140000 ;
    END

# P/G pin shape extracted from block 'tcam_32x28'
    PORT
      LAYER met4 ;
        RECT 1296.825000 2129.320000 1298.565000 2517.300000 ;
      LAYER met4 ;
        RECT 828.305000 2129.320000 830.045000 2517.300000 ;
      LAYER met3 ;
        RECT 828.305000 2129.320000 1298.565000 2131.060000 ;
      LAYER met3 ;
        RECT 828.305000 2515.560000 1298.565000 2517.300000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1858.965000 2129.415000 1860.705000 2517.395000 ;
      LAYER met4 ;
        RECT 1390.445000 2129.415000 1392.185000 2517.395000 ;
      LAYER met3 ;
        RECT 1390.445000 2129.415000 1860.705000 2131.155000 ;
      LAYER met3 ;
        RECT 1390.445000 2515.655000 1860.705000 2517.395000 ;
    END
    PORT
      LAYER met4 ;
        RECT 802.635000 2090.285000 804.635000 2552.525000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1884.575000 2090.285000 1886.575000 2552.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 802.635000 2550.525000 1886.575000 2552.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 802.635000 2090.285000 1886.575000 2092.285000 ;
    END
# end of P/G pin shape extracted from block 'tcam_32x28'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 1425.540000 472.830000 1895.800000 474.570000 ;
      LAYER met3 ;
        RECT 1425.540000 86.590000 1895.800000 88.330000 ;
      LAYER met4 ;
        RECT 1425.540000 86.590000 1427.280000 474.570000 ;
      LAYER met4 ;
        RECT 1894.060000 86.590000 1895.800000 474.570000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 1425.540000 982.530000 1895.800000 984.270000 ;
      LAYER met3 ;
        RECT 1425.540000 596.290000 1895.800000 598.030000 ;
      LAYER met4 ;
        RECT 1425.540000 596.290000 1427.280000 984.270000 ;
      LAYER met4 ;
        RECT 1894.060000 596.290000 1895.800000 984.270000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 1425.540000 1492.230000 1895.800000 1493.970000 ;
      LAYER met3 ;
        RECT 1425.540000 1105.990000 1895.800000 1107.730000 ;
      LAYER met4 ;
        RECT 1425.540000 1105.990000 1427.280000 1493.970000 ;
      LAYER met4 ;
        RECT 1894.060000 1105.990000 1895.800000 1493.970000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 1425.540000 2001.930000 1895.800000 2003.670000 ;
      LAYER met3 ;
        RECT 1425.540000 1615.690000 1895.800000 1617.430000 ;
      LAYER met4 ;
        RECT 1425.540000 1615.690000 1427.280000 2003.670000 ;
      LAYER met4 ;
        RECT 1894.060000 1615.690000 1895.800000 2003.670000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 792.760000 472.830000 1263.020000 474.570000 ;
      LAYER met3 ;
        RECT 792.760000 86.590000 1263.020000 88.330000 ;
      LAYER met4 ;
        RECT 792.760000 86.590000 794.500000 474.570000 ;
      LAYER met4 ;
        RECT 1261.280000 86.590000 1263.020000 474.570000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 792.760000 982.530000 1263.020000 984.270000 ;
      LAYER met3 ;
        RECT 792.760000 596.290000 1263.020000 598.030000 ;
      LAYER met4 ;
        RECT 792.760000 596.290000 794.500000 984.270000 ;
      LAYER met4 ;
        RECT 1261.280000 596.290000 1263.020000 984.270000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 792.760000 1492.230000 1263.020000 1493.970000 ;
      LAYER met3 ;
        RECT 792.760000 1105.990000 1263.020000 1107.730000 ;
      LAYER met4 ;
        RECT 792.760000 1105.990000 794.500000 1493.970000 ;
      LAYER met4 ;
        RECT 1261.280000 1105.990000 1263.020000 1493.970000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 792.760000 2001.930000 1263.020000 2003.670000 ;
      LAYER met3 ;
        RECT 792.760000 1615.690000 1263.020000 1617.430000 ;
      LAYER met4 ;
        RECT 792.760000 1615.690000 794.500000 2003.670000 ;
      LAYER met4 ;
        RECT 1261.280000 1615.690000 1263.020000 2003.670000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END vccd1
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 1926.480000 2595.220000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 1926.480000 2595.220000 ;
    LAYER met2 ;
      RECT 1921.310000 2594.595000 1926.480000 2595.220000 ;
      RECT 1869.410000 2594.595000 1920.890000 2595.220000 ;
      RECT 3.910000 2594.595000 54.690000 2595.220000 ;
      RECT 0.000000 2594.595000 3.490000 2595.220000 ;
      RECT 1869.410000 2594.590000 1926.480000 2594.595000 ;
      RECT 1814.510000 2594.590000 1868.990000 2595.220000 ;
      RECT 1759.510000 2594.590000 1814.090000 2595.220000 ;
      RECT 1704.510000 2594.590000 1759.090000 2595.220000 ;
      RECT 1649.410000 2594.590000 1704.090000 2595.220000 ;
      RECT 1594.510000 2594.590000 1648.990000 2595.220000 ;
      RECT 1539.510000 2594.590000 1594.090000 2595.220000 ;
      RECT 1484.510000 2594.590000 1539.090000 2595.220000 ;
      RECT 1429.510000 2594.590000 1484.090000 2595.220000 ;
      RECT 1374.610000 2594.590000 1429.090000 2595.220000 ;
      RECT 1319.610000 2594.590000 1374.190000 2595.220000 ;
      RECT 1264.610000 2594.590000 1319.190000 2595.220000 ;
      RECT 1209.610000 2594.590000 1264.190000 2595.220000 ;
      RECT 1154.710000 2594.590000 1209.190000 2595.220000 ;
      RECT 1099.710000 2594.590000 1154.290000 2595.220000 ;
      RECT 1044.710000 2594.590000 1099.290000 2595.220000 ;
      RECT 989.710000 2594.590000 1044.290000 2595.220000 ;
      RECT 934.810000 2594.590000 989.290000 2595.220000 ;
      RECT 879.810000 2594.590000 934.390000 2595.220000 ;
      RECT 824.810000 2594.590000 879.390000 2595.220000 ;
      RECT 769.710000 2594.590000 824.390000 2595.220000 ;
      RECT 714.710000 2594.590000 769.290000 2595.220000 ;
      RECT 659.810000 2594.590000 714.290000 2595.220000 ;
      RECT 604.810000 2594.590000 659.390000 2595.220000 ;
      RECT 549.810000 2594.590000 604.390000 2595.220000 ;
      RECT 494.810000 2594.590000 549.390000 2595.220000 ;
      RECT 439.910000 2594.590000 494.390000 2595.220000 ;
      RECT 384.910000 2594.590000 439.490000 2595.220000 ;
      RECT 329.910000 2594.590000 384.490000 2595.220000 ;
      RECT 274.910000 2594.590000 329.490000 2595.220000 ;
      RECT 220.010000 2594.590000 274.490000 2595.220000 ;
      RECT 165.010000 2594.590000 219.590000 2595.220000 ;
      RECT 110.010000 2594.590000 164.590000 2595.220000 ;
      RECT 55.110000 2594.590000 109.590000 2595.220000 ;
      RECT 0.000000 2594.590000 54.690000 2594.595000 ;
      RECT 0.000000 0.630000 1926.480000 2594.590000 ;
      RECT 1920.410000 0.625000 1926.480000 0.630000 ;
      RECT 0.000000 0.625000 3.590000 0.630000 ;
      RECT 1923.010000 0.000000 1926.480000 0.625000 ;
      RECT 1920.410000 0.000000 1922.590000 0.625000 ;
      RECT 1916.510000 0.000000 1919.990000 0.630000 ;
      RECT 1912.610000 0.000000 1916.090000 0.630000 ;
      RECT 1908.810000 0.000000 1912.190000 0.630000 ;
      RECT 1904.910000 0.000000 1908.390000 0.630000 ;
      RECT 1901.010000 0.000000 1904.490000 0.630000 ;
      RECT 1897.010000 0.000000 1900.590000 0.630000 ;
      RECT 1893.110000 0.000000 1896.590000 0.630000 ;
      RECT 1889.210000 0.000000 1892.690000 0.630000 ;
      RECT 1885.310000 0.000000 1888.790000 0.630000 ;
      RECT 1881.410000 0.000000 1884.890000 0.630000 ;
      RECT 1877.510000 0.000000 1880.990000 0.630000 ;
      RECT 1873.610000 0.000000 1877.090000 0.630000 ;
      RECT 1869.710000 0.000000 1873.190000 0.630000 ;
      RECT 1865.810000 0.000000 1869.290000 0.630000 ;
      RECT 1861.910000 0.000000 1865.390000 0.630000 ;
      RECT 1858.010000 0.000000 1861.490000 0.630000 ;
      RECT 1854.110000 0.000000 1857.590000 0.630000 ;
      RECT 1850.210000 0.000000 1853.690000 0.630000 ;
      RECT 1846.310000 0.000000 1849.790000 0.630000 ;
      RECT 1842.410000 0.000000 1845.890000 0.630000 ;
      RECT 1838.510000 0.000000 1841.990000 0.630000 ;
      RECT 1834.610000 0.000000 1838.090000 0.630000 ;
      RECT 1830.710000 0.000000 1834.190000 0.630000 ;
      RECT 1826.810000 0.000000 1830.290000 0.630000 ;
      RECT 1822.910000 0.000000 1826.390000 0.630000 ;
      RECT 1818.910000 0.000000 1822.490000 0.630000 ;
      RECT 1815.010000 0.000000 1818.490000 0.630000 ;
      RECT 1811.110000 0.000000 1814.590000 0.630000 ;
      RECT 1807.210000 0.000000 1810.690000 0.630000 ;
      RECT 1803.310000 0.000000 1806.790000 0.630000 ;
      RECT 1799.510000 0.000000 1802.890000 0.630000 ;
      RECT 1795.610000 0.000000 1799.090000 0.630000 ;
      RECT 1791.610000 0.000000 1795.190000 0.630000 ;
      RECT 1787.810000 0.000000 1791.190000 0.630000 ;
      RECT 1783.910000 0.000000 1787.390000 0.630000 ;
      RECT 1780.010000 0.000000 1783.490000 0.630000 ;
      RECT 1776.110000 0.000000 1779.590000 0.630000 ;
      RECT 1772.210000 0.000000 1775.690000 0.630000 ;
      RECT 1768.210000 0.000000 1771.790000 0.630000 ;
      RECT 1764.310000 0.000000 1767.790000 0.630000 ;
      RECT 1760.410000 0.000000 1763.890000 0.630000 ;
      RECT 1756.510000 0.000000 1759.990000 0.630000 ;
      RECT 1752.610000 0.000000 1756.090000 0.630000 ;
      RECT 1748.710000 0.000000 1752.190000 0.630000 ;
      RECT 1744.810000 0.000000 1748.290000 0.630000 ;
      RECT 1740.810000 0.000000 1744.390000 0.630000 ;
      RECT 1736.910000 0.000000 1740.390000 0.630000 ;
      RECT 1733.010000 0.000000 1736.490000 0.630000 ;
      RECT 1729.210000 0.000000 1732.590000 0.630000 ;
      RECT 1725.310000 0.000000 1728.790000 0.630000 ;
      RECT 1721.510000 0.000000 1724.890000 0.630000 ;
      RECT 1717.610000 0.000000 1721.090000 0.630000 ;
      RECT 1713.610000 0.000000 1717.190000 0.630000 ;
      RECT 1709.710000 0.000000 1713.190000 0.630000 ;
      RECT 1705.810000 0.000000 1709.290000 0.630000 ;
      RECT 1701.910000 0.000000 1705.390000 0.630000 ;
      RECT 1698.010000 0.000000 1701.490000 0.630000 ;
      RECT 1694.110000 0.000000 1697.590000 0.630000 ;
      RECT 1690.110000 0.000000 1693.690000 0.630000 ;
      RECT 1686.210000 0.000000 1689.690000 0.630000 ;
      RECT 1682.310000 0.000000 1685.790000 0.630000 ;
      RECT 1678.410000 0.000000 1681.890000 0.630000 ;
      RECT 1674.510000 0.000000 1677.990000 0.630000 ;
      RECT 1670.610000 0.000000 1674.090000 0.630000 ;
      RECT 1666.710000 0.000000 1670.190000 0.630000 ;
      RECT 1662.810000 0.000000 1666.290000 0.630000 ;
      RECT 1658.910000 0.000000 1662.390000 0.630000 ;
      RECT 1655.110000 0.000000 1658.490000 0.630000 ;
      RECT 1651.210000 0.000000 1654.690000 0.630000 ;
      RECT 1647.310000 0.000000 1650.790000 0.630000 ;
      RECT 1643.410000 0.000000 1646.890000 0.630000 ;
      RECT 1639.510000 0.000000 1642.990000 0.630000 ;
      RECT 1635.510000 0.000000 1639.090000 0.630000 ;
      RECT 1631.610000 0.000000 1635.090000 0.630000 ;
      RECT 1627.710000 0.000000 1631.190000 0.630000 ;
      RECT 1623.810000 0.000000 1627.290000 0.630000 ;
      RECT 1619.910000 0.000000 1623.390000 0.630000 ;
      RECT 1616.010000 0.000000 1619.490000 0.630000 ;
      RECT 1612.010000 0.000000 1615.590000 0.630000 ;
      RECT 1608.110000 0.000000 1611.590000 0.630000 ;
      RECT 1604.210000 0.000000 1607.690000 0.630000 ;
      RECT 1600.410000 0.000000 1603.790000 0.630000 ;
      RECT 1596.510000 0.000000 1599.990000 0.630000 ;
      RECT 1592.610000 0.000000 1596.090000 0.630000 ;
      RECT 1588.710000 0.000000 1592.190000 0.630000 ;
      RECT 1584.810000 0.000000 1588.290000 0.630000 ;
      RECT 1580.910000 0.000000 1584.390000 0.630000 ;
      RECT 1577.010000 0.000000 1580.490000 0.630000 ;
      RECT 1573.110000 0.000000 1576.590000 0.630000 ;
      RECT 1569.210000 0.000000 1572.690000 0.630000 ;
      RECT 1565.310000 0.000000 1568.790000 0.630000 ;
      RECT 1561.410000 0.000000 1564.890000 0.630000 ;
      RECT 1557.410000 0.000000 1560.990000 0.630000 ;
      RECT 1553.510000 0.000000 1556.990000 0.630000 ;
      RECT 1549.610000 0.000000 1553.090000 0.630000 ;
      RECT 1545.710000 0.000000 1549.190000 0.630000 ;
      RECT 1541.810000 0.000000 1545.290000 0.630000 ;
      RECT 1538.010000 0.000000 1541.390000 0.630000 ;
      RECT 1534.010000 0.000000 1537.590000 0.630000 ;
      RECT 1530.110000 0.000000 1533.590000 0.630000 ;
      RECT 1526.210000 0.000000 1529.690000 0.630000 ;
      RECT 1522.310000 0.000000 1525.790000 0.630000 ;
      RECT 1518.410000 0.000000 1521.890000 0.630000 ;
      RECT 1514.510000 0.000000 1517.990000 0.630000 ;
      RECT 1510.710000 0.000000 1514.090000 0.630000 ;
      RECT 1506.710000 0.000000 1510.290000 0.630000 ;
      RECT 1502.810000 0.000000 1506.290000 0.630000 ;
      RECT 1498.910000 0.000000 1502.390000 0.630000 ;
      RECT 1495.010000 0.000000 1498.490000 0.630000 ;
      RECT 1491.110000 0.000000 1494.590000 0.630000 ;
      RECT 1487.210000 0.000000 1490.690000 0.630000 ;
      RECT 1483.310000 0.000000 1486.790000 0.630000 ;
      RECT 1479.410000 0.000000 1482.890000 0.630000 ;
      RECT 1475.510000 0.000000 1478.990000 0.630000 ;
      RECT 1471.610000 0.000000 1475.090000 0.630000 ;
      RECT 1467.710000 0.000000 1471.190000 0.630000 ;
      RECT 1463.810000 0.000000 1467.290000 0.630000 ;
      RECT 1459.910000 0.000000 1463.390000 0.630000 ;
      RECT 1455.910000 0.000000 1459.490000 0.630000 ;
      RECT 1452.010000 0.000000 1455.490000 0.630000 ;
      RECT 1448.110000 0.000000 1451.590000 0.630000 ;
      RECT 1444.210000 0.000000 1447.690000 0.630000 ;
      RECT 1440.410000 0.000000 1443.790000 0.630000 ;
      RECT 1436.510000 0.000000 1439.990000 0.630000 ;
      RECT 1432.610000 0.000000 1436.090000 0.630000 ;
      RECT 1428.610000 0.000000 1432.190000 0.630000 ;
      RECT 1424.710000 0.000000 1428.190000 0.630000 ;
      RECT 1420.810000 0.000000 1424.290000 0.630000 ;
      RECT 1417.010000 0.000000 1420.390000 0.630000 ;
      RECT 1413.110000 0.000000 1416.590000 0.630000 ;
      RECT 1409.210000 0.000000 1412.690000 0.630000 ;
      RECT 1405.310000 0.000000 1408.790000 0.630000 ;
      RECT 1401.310000 0.000000 1404.890000 0.630000 ;
      RECT 1397.410000 0.000000 1400.890000 0.630000 ;
      RECT 1393.510000 0.000000 1396.990000 0.630000 ;
      RECT 1389.610000 0.000000 1393.090000 0.630000 ;
      RECT 1385.710000 0.000000 1389.190000 0.630000 ;
      RECT 1381.810000 0.000000 1385.290000 0.630000 ;
      RECT 1377.810000 0.000000 1381.390000 0.630000 ;
      RECT 1373.910000 0.000000 1377.390000 0.630000 ;
      RECT 1370.110000 0.000000 1373.490000 0.630000 ;
      RECT 1366.210000 0.000000 1369.690000 0.630000 ;
      RECT 1362.310000 0.000000 1365.790000 0.630000 ;
      RECT 1358.410000 0.000000 1361.890000 0.630000 ;
      RECT 1354.510000 0.000000 1357.990000 0.630000 ;
      RECT 1350.610000 0.000000 1354.090000 0.630000 ;
      RECT 1346.710000 0.000000 1350.190000 0.630000 ;
      RECT 1342.810000 0.000000 1346.290000 0.630000 ;
      RECT 1338.910000 0.000000 1342.390000 0.630000 ;
      RECT 1335.010000 0.000000 1338.490000 0.630000 ;
      RECT 1331.110000 0.000000 1334.590000 0.630000 ;
      RECT 1327.210000 0.000000 1330.690000 0.630000 ;
      RECT 1323.210000 0.000000 1326.790000 0.630000 ;
      RECT 1319.310000 0.000000 1322.790000 0.630000 ;
      RECT 1315.410000 0.000000 1318.890000 0.630000 ;
      RECT 1311.510000 0.000000 1314.990000 0.630000 ;
      RECT 1307.610000 0.000000 1311.090000 0.630000 ;
      RECT 1303.710000 0.000000 1307.190000 0.630000 ;
      RECT 1299.810000 0.000000 1303.290000 0.630000 ;
      RECT 1296.010000 0.000000 1299.390000 0.630000 ;
      RECT 1292.110000 0.000000 1295.590000 0.630000 ;
      RECT 1288.210000 0.000000 1291.690000 0.630000 ;
      RECT 1284.310000 0.000000 1287.790000 0.630000 ;
      RECT 1280.410000 0.000000 1283.890000 0.630000 ;
      RECT 1276.510000 0.000000 1279.990000 0.630000 ;
      RECT 1272.510000 0.000000 1276.090000 0.630000 ;
      RECT 1268.610000 0.000000 1272.090000 0.630000 ;
      RECT 1264.710000 0.000000 1268.190000 0.630000 ;
      RECT 1260.810000 0.000000 1264.290000 0.630000 ;
      RECT 1256.910000 0.000000 1260.390000 0.630000 ;
      RECT 1253.010000 0.000000 1256.490000 0.630000 ;
      RECT 1249.110000 0.000000 1252.590000 0.630000 ;
      RECT 1245.110000 0.000000 1248.690000 0.630000 ;
      RECT 1241.210000 0.000000 1244.690000 0.630000 ;
      RECT 1237.310000 0.000000 1240.790000 0.630000 ;
      RECT 1233.410000 0.000000 1236.890000 0.630000 ;
      RECT 1229.610000 0.000000 1232.990000 0.630000 ;
      RECT 1225.710000 0.000000 1229.190000 0.630000 ;
      RECT 1221.810000 0.000000 1225.290000 0.630000 ;
      RECT 1217.910000 0.000000 1221.390000 0.630000 ;
      RECT 1214.010000 0.000000 1217.490000 0.630000 ;
      RECT 1210.110000 0.000000 1213.590000 0.630000 ;
      RECT 1206.210000 0.000000 1209.690000 0.630000 ;
      RECT 1202.310000 0.000000 1205.790000 0.630000 ;
      RECT 1198.410000 0.000000 1201.890000 0.630000 ;
      RECT 1194.410000 0.000000 1197.990000 0.630000 ;
      RECT 1190.510000 0.000000 1193.990000 0.630000 ;
      RECT 1186.610000 0.000000 1190.090000 0.630000 ;
      RECT 1182.710000 0.000000 1186.190000 0.630000 ;
      RECT 1178.810000 0.000000 1182.290000 0.630000 ;
      RECT 1174.910000 0.000000 1178.390000 0.630000 ;
      RECT 1171.010000 0.000000 1174.490000 0.630000 ;
      RECT 1167.110000 0.000000 1170.590000 0.630000 ;
      RECT 1163.210000 0.000000 1166.690000 0.630000 ;
      RECT 1159.310000 0.000000 1162.790000 0.630000 ;
      RECT 1155.410000 0.000000 1158.890000 0.630000 ;
      RECT 1151.610000 0.000000 1154.990000 0.630000 ;
      RECT 1147.710000 0.000000 1151.190000 0.630000 ;
      RECT 1143.710000 0.000000 1147.290000 0.630000 ;
      RECT 1139.810000 0.000000 1143.290000 0.630000 ;
      RECT 1135.910000 0.000000 1139.390000 0.630000 ;
      RECT 1132.010000 0.000000 1135.490000 0.630000 ;
      RECT 1128.110000 0.000000 1131.590000 0.630000 ;
      RECT 1124.210000 0.000000 1127.690000 0.630000 ;
      RECT 1120.310000 0.000000 1123.790000 0.630000 ;
      RECT 1116.310000 0.000000 1119.890000 0.630000 ;
      RECT 1112.410000 0.000000 1115.890000 0.630000 ;
      RECT 1108.610000 0.000000 1111.990000 0.630000 ;
      RECT 1104.710000 0.000000 1108.190000 0.630000 ;
      RECT 1100.810000 0.000000 1104.290000 0.630000 ;
      RECT 1096.910000 0.000000 1100.390000 0.630000 ;
      RECT 1093.010000 0.000000 1096.490000 0.630000 ;
      RECT 1089.010000 0.000000 1092.590000 0.630000 ;
      RECT 1085.110000 0.000000 1088.590000 0.630000 ;
      RECT 1081.310000 0.000000 1084.690000 0.630000 ;
      RECT 1077.410000 0.000000 1080.890000 0.630000 ;
      RECT 1073.510000 0.000000 1076.990000 0.630000 ;
      RECT 1069.610000 0.000000 1073.090000 0.630000 ;
      RECT 1065.610000 0.000000 1069.190000 0.630000 ;
      RECT 1061.710000 0.000000 1065.190000 0.630000 ;
      RECT 1057.810000 0.000000 1061.290000 0.630000 ;
      RECT 1053.910000 0.000000 1057.390000 0.630000 ;
      RECT 1050.010000 0.000000 1053.490000 0.630000 ;
      RECT 1046.210000 0.000000 1049.590000 0.630000 ;
      RECT 1042.310000 0.000000 1045.790000 0.630000 ;
      RECT 1038.310000 0.000000 1041.890000 0.630000 ;
      RECT 1034.410000 0.000000 1037.890000 0.630000 ;
      RECT 1030.510000 0.000000 1033.990000 0.630000 ;
      RECT 1026.610000 0.000000 1030.090000 0.630000 ;
      RECT 1022.710000 0.000000 1026.190000 0.630000 ;
      RECT 1018.810000 0.000000 1022.290000 0.630000 ;
      RECT 1014.910000 0.000000 1018.390000 0.630000 ;
      RECT 1011.010000 0.000000 1014.490000 0.630000 ;
      RECT 1007.110000 0.000000 1010.590000 0.630000 ;
      RECT 1003.210000 0.000000 1006.690000 0.630000 ;
      RECT 999.310000 0.000000 1002.790000 0.630000 ;
      RECT 995.410000 0.000000 998.890000 0.630000 ;
      RECT 991.510000 0.000000 994.990000 0.630000 ;
      RECT 987.610000 0.000000 991.090000 0.630000 ;
      RECT 983.710000 0.000000 987.190000 0.630000 ;
      RECT 979.810000 0.000000 983.290000 0.630000 ;
      RECT 975.910000 0.000000 979.390000 0.630000 ;
      RECT 972.010000 0.000000 975.490000 0.630000 ;
      RECT 968.110000 0.000000 971.590000 0.630000 ;
      RECT 964.210000 0.000000 967.690000 0.630000 ;
      RECT 960.210000 0.000000 963.790000 0.630000 ;
      RECT 956.310000 0.000000 959.790000 0.630000 ;
      RECT 952.410000 0.000000 955.890000 0.630000 ;
      RECT 948.510000 0.000000 951.990000 0.630000 ;
      RECT 944.610000 0.000000 948.090000 0.630000 ;
      RECT 940.710000 0.000000 944.190000 0.630000 ;
      RECT 936.910000 0.000000 940.290000 0.630000 ;
      RECT 932.910000 0.000000 936.490000 0.630000 ;
      RECT 929.010000 0.000000 932.490000 0.630000 ;
      RECT 925.210000 0.000000 928.590000 0.630000 ;
      RECT 921.310000 0.000000 924.790000 0.630000 ;
      RECT 917.410000 0.000000 920.890000 0.630000 ;
      RECT 913.510000 0.000000 916.990000 0.630000 ;
      RECT 909.510000 0.000000 913.090000 0.630000 ;
      RECT 905.610000 0.000000 909.090000 0.630000 ;
      RECT 901.710000 0.000000 905.190000 0.630000 ;
      RECT 897.810000 0.000000 901.290000 0.630000 ;
      RECT 893.910000 0.000000 897.390000 0.630000 ;
      RECT 890.010000 0.000000 893.490000 0.630000 ;
      RECT 886.110000 0.000000 889.590000 0.630000 ;
      RECT 882.110000 0.000000 885.690000 0.630000 ;
      RECT 878.210000 0.000000 881.690000 0.630000 ;
      RECT 874.310000 0.000000 877.790000 0.630000 ;
      RECT 870.410000 0.000000 873.890000 0.630000 ;
      RECT 866.610000 0.000000 869.990000 0.630000 ;
      RECT 862.810000 0.000000 866.190000 0.630000 ;
      RECT 858.910000 0.000000 862.390000 0.630000 ;
      RECT 854.910000 0.000000 858.490000 0.630000 ;
      RECT 851.010000 0.000000 854.490000 0.630000 ;
      RECT 847.110000 0.000000 850.590000 0.630000 ;
      RECT 843.210000 0.000000 846.690000 0.630000 ;
      RECT 839.310000 0.000000 842.790000 0.630000 ;
      RECT 835.410000 0.000000 838.890000 0.630000 ;
      RECT 831.410000 0.000000 834.990000 0.630000 ;
      RECT 827.510000 0.000000 830.990000 0.630000 ;
      RECT 823.610000 0.000000 827.090000 0.630000 ;
      RECT 819.710000 0.000000 823.190000 0.630000 ;
      RECT 815.810000 0.000000 819.290000 0.630000 ;
      RECT 811.910000 0.000000 815.390000 0.630000 ;
      RECT 808.010000 0.000000 811.490000 0.630000 ;
      RECT 804.110000 0.000000 807.590000 0.630000 ;
      RECT 800.210000 0.000000 803.690000 0.630000 ;
      RECT 796.310000 0.000000 799.790000 0.630000 ;
      RECT 792.510000 0.000000 795.890000 0.630000 ;
      RECT 788.610000 0.000000 792.090000 0.630000 ;
      RECT 784.710000 0.000000 788.190000 0.630000 ;
      RECT 780.810000 0.000000 784.290000 0.630000 ;
      RECT 776.810000 0.000000 780.390000 0.630000 ;
      RECT 772.910000 0.000000 776.390000 0.630000 ;
      RECT 769.010000 0.000000 772.490000 0.630000 ;
      RECT 765.110000 0.000000 768.590000 0.630000 ;
      RECT 761.210000 0.000000 764.690000 0.630000 ;
      RECT 757.310000 0.000000 760.790000 0.630000 ;
      RECT 753.310000 0.000000 756.890000 0.630000 ;
      RECT 749.410000 0.000000 752.890000 0.630000 ;
      RECT 745.510000 0.000000 748.990000 0.630000 ;
      RECT 741.710000 0.000000 745.090000 0.630000 ;
      RECT 737.810000 0.000000 741.290000 0.630000 ;
      RECT 733.910000 0.000000 737.390000 0.630000 ;
      RECT 730.010000 0.000000 733.490000 0.630000 ;
      RECT 726.010000 0.000000 729.590000 0.630000 ;
      RECT 722.210000 0.000000 725.590000 0.630000 ;
      RECT 718.310000 0.000000 721.790000 0.630000 ;
      RECT 714.410000 0.000000 717.890000 0.630000 ;
      RECT 710.510000 0.000000 713.990000 0.630000 ;
      RECT 706.610000 0.000000 710.090000 0.630000 ;
      RECT 702.710000 0.000000 706.190000 0.630000 ;
      RECT 698.710000 0.000000 702.290000 0.630000 ;
      RECT 694.810000 0.000000 698.290000 0.630000 ;
      RECT 690.910000 0.000000 694.390000 0.630000 ;
      RECT 687.010000 0.000000 690.490000 0.630000 ;
      RECT 683.110000 0.000000 686.590000 0.630000 ;
      RECT 679.210000 0.000000 682.690000 0.630000 ;
      RECT 675.310000 0.000000 678.790000 0.630000 ;
      RECT 671.410000 0.000000 674.890000 0.630000 ;
      RECT 667.510000 0.000000 670.990000 0.630000 ;
      RECT 663.610000 0.000000 667.090000 0.630000 ;
      RECT 659.710000 0.000000 663.190000 0.630000 ;
      RECT 655.810000 0.000000 659.290000 0.630000 ;
      RECT 651.910000 0.000000 655.390000 0.630000 ;
      RECT 648.010000 0.000000 651.490000 0.630000 ;
      RECT 644.110000 0.000000 647.590000 0.630000 ;
      RECT 640.210000 0.000000 643.690000 0.630000 ;
      RECT 636.310000 0.000000 639.790000 0.630000 ;
      RECT 632.410000 0.000000 635.890000 0.630000 ;
      RECT 628.510000 0.000000 631.990000 0.630000 ;
      RECT 624.610000 0.000000 628.090000 0.630000 ;
      RECT 620.710000 0.000000 624.190000 0.630000 ;
      RECT 616.810000 0.000000 620.290000 0.630000 ;
      RECT 612.910000 0.000000 616.390000 0.630000 ;
      RECT 609.010000 0.000000 612.490000 0.630000 ;
      RECT 605.110000 0.000000 608.590000 0.630000 ;
      RECT 601.210000 0.000000 604.690000 0.630000 ;
      RECT 597.210000 0.000000 600.790000 0.630000 ;
      RECT 593.310000 0.000000 596.790000 0.630000 ;
      RECT 589.410000 0.000000 592.890000 0.630000 ;
      RECT 585.510000 0.000000 588.990000 0.630000 ;
      RECT 581.610000 0.000000 585.090000 0.630000 ;
      RECT 577.810000 0.000000 581.190000 0.630000 ;
      RECT 573.910000 0.000000 577.390000 0.630000 ;
      RECT 569.910000 0.000000 573.490000 0.630000 ;
      RECT 566.010000 0.000000 569.490000 0.630000 ;
      RECT 562.110000 0.000000 565.590000 0.630000 ;
      RECT 558.210000 0.000000 561.690000 0.630000 ;
      RECT 554.410000 0.000000 557.790000 0.630000 ;
      RECT 550.510000 0.000000 553.990000 0.630000 ;
      RECT 546.610000 0.000000 550.090000 0.630000 ;
      RECT 542.610000 0.000000 546.190000 0.630000 ;
      RECT 538.710000 0.000000 542.190000 0.630000 ;
      RECT 534.810000 0.000000 538.290000 0.630000 ;
      RECT 530.910000 0.000000 534.390000 0.630000 ;
      RECT 527.010000 0.000000 530.490000 0.630000 ;
      RECT 523.110000 0.000000 526.590000 0.630000 ;
      RECT 519.110000 0.000000 522.690000 0.630000 ;
      RECT 515.210000 0.000000 518.690000 0.630000 ;
      RECT 511.310000 0.000000 514.790000 0.630000 ;
      RECT 507.510000 0.000000 510.890000 0.630000 ;
      RECT 503.610000 0.000000 507.090000 0.630000 ;
      RECT 499.710000 0.000000 503.190000 0.630000 ;
      RECT 495.810000 0.000000 499.290000 0.630000 ;
      RECT 491.910000 0.000000 495.390000 0.630000 ;
      RECT 488.010000 0.000000 491.490000 0.630000 ;
      RECT 484.110000 0.000000 487.590000 0.630000 ;
      RECT 480.210000 0.000000 483.690000 0.630000 ;
      RECT 476.310000 0.000000 479.790000 0.630000 ;
      RECT 472.410000 0.000000 475.890000 0.630000 ;
      RECT 468.510000 0.000000 471.990000 0.630000 ;
      RECT 464.510000 0.000000 468.090000 0.630000 ;
      RECT 460.610000 0.000000 464.090000 0.630000 ;
      RECT 456.710000 0.000000 460.190000 0.630000 ;
      RECT 452.810000 0.000000 456.290000 0.630000 ;
      RECT 448.910000 0.000000 452.390000 0.630000 ;
      RECT 445.010000 0.000000 448.490000 0.630000 ;
      RECT 441.010000 0.000000 444.590000 0.630000 ;
      RECT 437.210000 0.000000 440.590000 0.630000 ;
      RECT 433.410000 0.000000 436.790000 0.630000 ;
      RECT 429.510000 0.000000 432.990000 0.630000 ;
      RECT 425.610000 0.000000 429.090000 0.630000 ;
      RECT 421.710000 0.000000 425.190000 0.630000 ;
      RECT 417.810000 0.000000 421.290000 0.630000 ;
      RECT 413.810000 0.000000 417.390000 0.630000 ;
      RECT 409.910000 0.000000 413.390000 0.630000 ;
      RECT 406.010000 0.000000 409.490000 0.630000 ;
      RECT 402.110000 0.000000 405.590000 0.630000 ;
      RECT 398.210000 0.000000 401.690000 0.630000 ;
      RECT 394.310000 0.000000 397.790000 0.630000 ;
      RECT 390.410000 0.000000 393.890000 0.630000 ;
      RECT 386.410000 0.000000 389.990000 0.630000 ;
      RECT 382.510000 0.000000 385.990000 0.630000 ;
      RECT 378.610000 0.000000 382.090000 0.630000 ;
      RECT 374.710000 0.000000 378.190000 0.630000 ;
      RECT 370.910000 0.000000 374.290000 0.630000 ;
      RECT 367.010000 0.000000 370.490000 0.630000 ;
      RECT 363.110000 0.000000 366.590000 0.630000 ;
      RECT 359.210000 0.000000 362.690000 0.630000 ;
      RECT 355.310000 0.000000 358.790000 0.630000 ;
      RECT 351.410000 0.000000 354.890000 0.630000 ;
      RECT 347.510000 0.000000 350.990000 0.630000 ;
      RECT 343.610000 0.000000 347.090000 0.630000 ;
      RECT 339.710000 0.000000 343.190000 0.630000 ;
      RECT 335.710000 0.000000 339.290000 0.630000 ;
      RECT 331.810000 0.000000 335.290000 0.630000 ;
      RECT 327.910000 0.000000 331.390000 0.630000 ;
      RECT 324.010000 0.000000 327.490000 0.630000 ;
      RECT 320.110000 0.000000 323.590000 0.630000 ;
      RECT 316.210000 0.000000 319.690000 0.630000 ;
      RECT 312.310000 0.000000 315.790000 0.630000 ;
      RECT 308.410000 0.000000 311.890000 0.630000 ;
      RECT 304.510000 0.000000 307.990000 0.630000 ;
      RECT 300.610000 0.000000 304.090000 0.630000 ;
      RECT 296.710000 0.000000 300.190000 0.630000 ;
      RECT 292.810000 0.000000 296.290000 0.630000 ;
      RECT 289.010000 0.000000 292.390000 0.630000 ;
      RECT 285.010000 0.000000 288.590000 0.630000 ;
      RECT 281.110000 0.000000 284.590000 0.630000 ;
      RECT 277.210000 0.000000 280.690000 0.630000 ;
      RECT 273.310000 0.000000 276.790000 0.630000 ;
      RECT 269.410000 0.000000 272.890000 0.630000 ;
      RECT 265.510000 0.000000 268.990000 0.630000 ;
      RECT 261.610000 0.000000 265.090000 0.630000 ;
      RECT 257.610000 0.000000 261.190000 0.630000 ;
      RECT 253.710000 0.000000 257.190000 0.630000 ;
      RECT 249.910000 0.000000 253.290000 0.630000 ;
      RECT 246.010000 0.000000 249.490000 0.630000 ;
      RECT 242.110000 0.000000 245.590000 0.630000 ;
      RECT 238.210000 0.000000 241.690000 0.630000 ;
      RECT 234.310000 0.000000 237.790000 0.630000 ;
      RECT 230.310000 0.000000 233.890000 0.630000 ;
      RECT 226.410000 0.000000 229.890000 0.630000 ;
      RECT 222.510000 0.000000 225.990000 0.630000 ;
      RECT 218.710000 0.000000 222.090000 0.630000 ;
      RECT 214.810000 0.000000 218.290000 0.630000 ;
      RECT 210.910000 0.000000 214.390000 0.630000 ;
      RECT 206.910000 0.000000 210.490000 0.630000 ;
      RECT 203.010000 0.000000 206.490000 0.630000 ;
      RECT 199.110000 0.000000 202.590000 0.630000 ;
      RECT 195.210000 0.000000 198.690000 0.630000 ;
      RECT 191.310000 0.000000 194.790000 0.630000 ;
      RECT 187.410000 0.000000 190.890000 0.630000 ;
      RECT 183.610000 0.000000 186.990000 0.630000 ;
      RECT 179.610000 0.000000 183.190000 0.630000 ;
      RECT 175.710000 0.000000 179.190000 0.630000 ;
      RECT 171.810000 0.000000 175.290000 0.630000 ;
      RECT 167.910000 0.000000 171.390000 0.630000 ;
      RECT 164.010000 0.000000 167.490000 0.630000 ;
      RECT 160.110000 0.000000 163.590000 0.630000 ;
      RECT 156.210000 0.000000 159.690000 0.630000 ;
      RECT 152.210000 0.000000 155.790000 0.630000 ;
      RECT 148.410000 0.000000 151.790000 0.630000 ;
      RECT 144.510000 0.000000 147.990000 0.630000 ;
      RECT 140.610000 0.000000 144.090000 0.630000 ;
      RECT 136.710000 0.000000 140.190000 0.630000 ;
      RECT 132.810000 0.000000 136.290000 0.630000 ;
      RECT 128.910000 0.000000 132.390000 0.630000 ;
      RECT 125.010000 0.000000 128.490000 0.630000 ;
      RECT 121.110000 0.000000 124.590000 0.630000 ;
      RECT 117.210000 0.000000 120.690000 0.630000 ;
      RECT 113.310000 0.000000 116.790000 0.630000 ;
      RECT 109.410000 0.000000 112.890000 0.630000 ;
      RECT 105.510000 0.000000 108.990000 0.630000 ;
      RECT 101.510000 0.000000 105.090000 0.630000 ;
      RECT 97.610000 0.000000 101.090000 0.630000 ;
      RECT 93.710000 0.000000 97.190000 0.630000 ;
      RECT 89.810000 0.000000 93.290000 0.630000 ;
      RECT 85.910000 0.000000 89.390000 0.630000 ;
      RECT 82.010000 0.000000 85.490000 0.630000 ;
      RECT 78.110000 0.000000 81.590000 0.630000 ;
      RECT 74.210000 0.000000 77.690000 0.630000 ;
      RECT 70.310000 0.000000 73.790000 0.630000 ;
      RECT 66.410000 0.000000 69.890000 0.630000 ;
      RECT 62.610000 0.000000 65.990000 0.630000 ;
      RECT 58.710000 0.000000 62.190000 0.630000 ;
      RECT 54.810000 0.000000 58.290000 0.630000 ;
      RECT 50.810000 0.000000 54.390000 0.630000 ;
      RECT 46.910000 0.000000 50.390000 0.630000 ;
      RECT 43.010000 0.000000 46.490000 0.630000 ;
      RECT 39.110000 0.000000 42.590000 0.630000 ;
      RECT 35.210000 0.000000 38.690000 0.630000 ;
      RECT 31.310000 0.000000 34.790000 0.630000 ;
      RECT 27.410000 0.000000 30.890000 0.630000 ;
      RECT 23.410000 0.000000 26.990000 0.630000 ;
      RECT 19.510000 0.000000 22.990000 0.630000 ;
      RECT 15.610000 0.000000 19.090000 0.630000 ;
      RECT 11.710000 0.000000 15.190000 0.630000 ;
      RECT 7.810000 0.000000 11.290000 0.630000 ;
      RECT 4.010000 0.000000 7.390000 0.630000 ;
      RECT 2.210000 0.000000 3.590000 0.625000 ;
      RECT 0.000000 0.000000 1.790000 0.625000 ;
    LAYER met3 ;
      RECT 0.000000 2587.340000 1926.480000 2595.220000 ;
      RECT 1919.900000 2582.540000 1926.480000 2587.340000 ;
      RECT 0.000000 2582.540000 6.580000 2587.340000 ;
      RECT 0.000000 2581.540000 1926.480000 2582.540000 ;
      RECT 1914.100000 2576.740000 1926.480000 2581.540000 ;
      RECT 0.000000 2576.740000 12.380000 2581.540000 ;
      RECT 0.000000 2524.000000 1926.480000 2576.740000 ;
      RECT 0.000000 2523.425000 1925.380000 2524.000000 ;
      RECT 1.100000 2523.100000 1925.380000 2523.425000 ;
      RECT 1.100000 2522.525000 1926.480000 2523.100000 ;
      RECT 0.000000 2478.305000 1926.480000 2522.525000 ;
      RECT 1.100000 2477.440000 1926.480000 2478.305000 ;
      RECT 1.100000 2477.405000 1925.380000 2477.440000 ;
      RECT 0.000000 2476.540000 1925.380000 2477.405000 ;
      RECT 0.000000 2430.785000 1926.480000 2476.540000 ;
      RECT 1.100000 2429.885000 1926.480000 2430.785000 ;
      RECT 0.000000 2428.865000 1926.480000 2429.885000 ;
      RECT 0.000000 2427.965000 1925.380000 2428.865000 ;
      RECT 0.000000 2383.075000 1926.480000 2427.965000 ;
      RECT 1.100000 2382.175000 1926.480000 2383.075000 ;
      RECT 0.000000 2380.385000 1926.480000 2382.175000 ;
      RECT 0.000000 2379.485000 1925.380000 2380.385000 ;
      RECT 0.000000 2335.265000 1926.480000 2379.485000 ;
      RECT 1.100000 2334.365000 1926.480000 2335.265000 ;
      RECT 0.000000 2331.715000 1926.480000 2334.365000 ;
      RECT 0.000000 2330.815000 1925.380000 2331.715000 ;
      RECT 0.000000 2287.745000 1926.480000 2330.815000 ;
      RECT 1.100000 2286.845000 1926.480000 2287.745000 ;
      RECT 0.000000 2283.040000 1926.480000 2286.845000 ;
      RECT 0.000000 2282.140000 1925.380000 2283.040000 ;
      RECT 0.000000 2240.035000 1926.480000 2282.140000 ;
      RECT 1.100000 2239.135000 1926.480000 2240.035000 ;
      RECT 0.000000 2234.465000 1926.480000 2239.135000 ;
      RECT 0.000000 2233.565000 1925.380000 2234.465000 ;
      RECT 0.000000 2192.420000 1926.480000 2233.565000 ;
      RECT 1.100000 2191.520000 1926.480000 2192.420000 ;
      RECT 0.000000 2185.985000 1926.480000 2191.520000 ;
      RECT 0.000000 2185.085000 1925.380000 2185.985000 ;
      RECT 0.000000 2144.705000 1926.480000 2185.085000 ;
      RECT 1.100000 2143.805000 1926.480000 2144.705000 ;
      RECT 0.000000 2137.410000 1926.480000 2143.805000 ;
      RECT 0.000000 2136.510000 1925.380000 2137.410000 ;
      RECT 0.000000 2097.090000 1926.480000 2136.510000 ;
      RECT 1.100000 2096.190000 1926.480000 2097.090000 ;
      RECT 0.000000 2088.740000 1926.480000 2096.190000 ;
      RECT 0.000000 2087.840000 1925.380000 2088.740000 ;
      RECT 0.000000 2049.280000 1926.480000 2087.840000 ;
      RECT 1.100000 2048.380000 1926.480000 2049.280000 ;
      RECT 0.000000 2040.260000 1926.480000 2048.380000 ;
      RECT 0.000000 2039.360000 1925.380000 2040.260000 ;
      RECT 0.000000 2001.760000 1926.480000 2039.360000 ;
      RECT 1.100000 2000.860000 1926.480000 2001.760000 ;
      RECT 0.000000 1991.680000 1926.480000 2000.860000 ;
      RECT 0.000000 1990.780000 1925.380000 1991.680000 ;
      RECT 0.000000 1954.050000 1926.480000 1990.780000 ;
      RECT 1.100000 1953.150000 1926.480000 1954.050000 ;
      RECT 0.000000 1943.105000 1926.480000 1953.150000 ;
      RECT 0.000000 1942.205000 1925.380000 1943.105000 ;
      RECT 0.000000 1906.435000 1926.480000 1942.205000 ;
      RECT 1.100000 1905.535000 1926.480000 1906.435000 ;
      RECT 0.000000 1894.720000 1926.480000 1905.535000 ;
      RECT 0.000000 1893.820000 1925.380000 1894.720000 ;
      RECT 0.000000 1858.820000 1926.480000 1893.820000 ;
      RECT 1.100000 1857.920000 1926.480000 1858.820000 ;
      RECT 0.000000 1845.955000 1926.480000 1857.920000 ;
      RECT 0.000000 1845.055000 1925.380000 1845.955000 ;
      RECT 0.000000 1811.105000 1926.480000 1845.055000 ;
      RECT 1.100000 1810.205000 1926.480000 1811.105000 ;
      RECT 0.000000 1797.380000 1926.480000 1810.205000 ;
      RECT 0.000000 1796.480000 1925.380000 1797.380000 ;
      RECT 0.000000 1763.490000 1926.480000 1796.480000 ;
      RECT 1.100000 1762.590000 1926.480000 1763.490000 ;
      RECT 0.000000 1748.800000 1926.480000 1762.590000 ;
      RECT 0.000000 1747.900000 1925.380000 1748.800000 ;
      RECT 0.000000 1715.780000 1926.480000 1747.900000 ;
      RECT 1.100000 1714.880000 1926.480000 1715.780000 ;
      RECT 0.000000 1700.320000 1926.480000 1714.880000 ;
      RECT 0.000000 1699.420000 1925.380000 1700.320000 ;
      RECT 0.000000 1668.260000 1926.480000 1699.420000 ;
      RECT 1.100000 1667.360000 1926.480000 1668.260000 ;
      RECT 0.000000 1651.650000 1926.480000 1667.360000 ;
      RECT 0.000000 1650.750000 1925.380000 1651.650000 ;
      RECT 0.000000 1620.545000 1926.480000 1650.750000 ;
      RECT 1.100000 1619.645000 1926.480000 1620.545000 ;
      RECT 0.000000 1602.980000 1926.480000 1619.645000 ;
      RECT 0.000000 1602.080000 1925.380000 1602.980000 ;
      RECT 0.000000 1572.930000 1926.480000 1602.080000 ;
      RECT 1.100000 1572.030000 1926.480000 1572.930000 ;
      RECT 0.000000 1554.595000 1926.480000 1572.030000 ;
      RECT 0.000000 1553.695000 1925.380000 1554.595000 ;
      RECT 0.000000 1525.120000 1926.480000 1553.695000 ;
      RECT 1.100000 1524.220000 1926.480000 1525.120000 ;
      RECT 0.000000 1505.920000 1926.480000 1524.220000 ;
      RECT 0.000000 1505.020000 1925.380000 1505.920000 ;
      RECT 0.000000 1477.410000 1926.480000 1505.020000 ;
      RECT 1.100000 1476.510000 1926.480000 1477.410000 ;
      RECT 0.000000 1457.440000 1926.480000 1476.510000 ;
      RECT 0.000000 1456.540000 1925.380000 1457.440000 ;
      RECT 0.000000 1429.795000 1926.480000 1456.540000 ;
      RECT 1.100000 1428.895000 1926.480000 1429.795000 ;
      RECT 0.000000 1408.675000 1926.480000 1428.895000 ;
      RECT 0.000000 1407.775000 1925.380000 1408.675000 ;
      RECT 0.000000 1382.180000 1926.480000 1407.775000 ;
      RECT 1.100000 1381.280000 1926.480000 1382.180000 ;
      RECT 0.000000 1360.290000 1926.480000 1381.280000 ;
      RECT 0.000000 1359.390000 1925.380000 1360.290000 ;
      RECT 0.000000 1334.465000 1926.480000 1359.390000 ;
      RECT 1.100000 1333.565000 1926.480000 1334.465000 ;
      RECT 0.000000 1311.620000 1926.480000 1333.565000 ;
      RECT 0.000000 1310.720000 1925.380000 1311.620000 ;
      RECT 0.000000 1286.850000 1926.480000 1310.720000 ;
      RECT 1.100000 1285.950000 1926.480000 1286.850000 ;
      RECT 0.000000 1263.040000 1926.480000 1285.950000 ;
      RECT 0.000000 1262.140000 1925.380000 1263.040000 ;
      RECT 0.000000 1239.330000 1926.480000 1262.140000 ;
      RECT 1.100000 1238.430000 1926.480000 1239.330000 ;
      RECT 0.000000 1214.660000 1926.480000 1238.430000 ;
      RECT 0.000000 1213.760000 1925.380000 1214.660000 ;
      RECT 0.000000 1191.620000 1926.480000 1213.760000 ;
      RECT 1.100000 1190.720000 1926.480000 1191.620000 ;
      RECT 0.000000 1165.985000 1926.480000 1190.720000 ;
      RECT 0.000000 1165.085000 1925.380000 1165.985000 ;
      RECT 0.000000 1144.100000 1926.480000 1165.085000 ;
      RECT 1.100000 1143.200000 1926.480000 1144.100000 ;
      RECT 0.000000 1117.315000 1926.480000 1143.200000 ;
      RECT 0.000000 1116.415000 1925.380000 1117.315000 ;
      RECT 0.000000 1096.385000 1926.480000 1116.415000 ;
      RECT 1.100000 1095.485000 1926.480000 1096.385000 ;
      RECT 0.000000 1068.740000 1926.480000 1095.485000 ;
      RECT 0.000000 1067.840000 1925.380000 1068.740000 ;
      RECT 0.000000 1048.580000 1926.480000 1067.840000 ;
      RECT 1.100000 1047.680000 1926.480000 1048.580000 ;
      RECT 0.000000 1020.260000 1926.480000 1047.680000 ;
      RECT 0.000000 1019.360000 1925.380000 1020.260000 ;
      RECT 0.000000 1000.865000 1926.480000 1019.360000 ;
      RECT 1.100000 999.965000 1926.480000 1000.865000 ;
      RECT 0.000000 971.585000 1926.480000 999.965000 ;
      RECT 0.000000 970.685000 1925.380000 971.585000 ;
      RECT 0.000000 953.250000 1926.480000 970.685000 ;
      RECT 1.100000 952.350000 1926.480000 953.250000 ;
      RECT 0.000000 923.010000 1926.480000 952.350000 ;
      RECT 0.000000 922.110000 1925.380000 923.010000 ;
      RECT 0.000000 905.540000 1926.480000 922.110000 ;
      RECT 1.100000 904.640000 1926.480000 905.540000 ;
      RECT 0.000000 874.530000 1926.480000 904.640000 ;
      RECT 0.000000 873.630000 1925.380000 874.530000 ;
      RECT 0.000000 857.920000 1926.480000 873.630000 ;
      RECT 1.100000 857.020000 1926.480000 857.920000 ;
      RECT 0.000000 825.955000 1926.480000 857.020000 ;
      RECT 0.000000 825.055000 1925.380000 825.955000 ;
      RECT 0.000000 810.210000 1926.480000 825.055000 ;
      RECT 1.100000 809.310000 1926.480000 810.210000 ;
      RECT 0.000000 777.280000 1926.480000 809.310000 ;
      RECT 0.000000 776.380000 1925.380000 777.280000 ;
      RECT 0.000000 762.595000 1926.480000 776.380000 ;
      RECT 1.100000 761.695000 1926.480000 762.595000 ;
      RECT 0.000000 728.900000 1926.480000 761.695000 ;
      RECT 0.000000 728.000000 1925.380000 728.900000 ;
      RECT 0.000000 715.075000 1926.480000 728.000000 ;
      RECT 1.100000 714.175000 1926.480000 715.075000 ;
      RECT 0.000000 680.225000 1926.480000 714.175000 ;
      RECT 0.000000 679.325000 1925.380000 680.225000 ;
      RECT 0.000000 667.460000 1926.480000 679.325000 ;
      RECT 1.100000 666.560000 1926.480000 667.460000 ;
      RECT 0.000000 631.650000 1926.480000 666.560000 ;
      RECT 0.000000 630.750000 1925.380000 631.650000 ;
      RECT 0.000000 619.745000 1926.480000 630.750000 ;
      RECT 1.100000 618.845000 1926.480000 619.745000 ;
      RECT 0.000000 583.075000 1926.480000 618.845000 ;
      RECT 0.000000 582.175000 1925.380000 583.075000 ;
      RECT 0.000000 572.130000 1926.480000 582.175000 ;
      RECT 1.100000 571.230000 1926.480000 572.130000 ;
      RECT 0.000000 534.500000 1926.480000 571.230000 ;
      RECT 0.000000 533.600000 1925.380000 534.500000 ;
      RECT 0.000000 524.420000 1926.480000 533.600000 ;
      RECT 1.100000 523.520000 1926.480000 524.420000 ;
      RECT 0.000000 485.825000 1926.480000 523.520000 ;
      RECT 0.000000 484.925000 1925.380000 485.825000 ;
      RECT 0.000000 476.610000 1926.480000 484.925000 ;
      RECT 1.100000 475.710000 1926.480000 476.610000 ;
      RECT 0.000000 437.345000 1926.480000 475.710000 ;
      RECT 0.000000 436.445000 1925.380000 437.345000 ;
      RECT 0.000000 429.090000 1926.480000 436.445000 ;
      RECT 1.100000 428.190000 1926.480000 429.090000 ;
      RECT 0.000000 388.675000 1926.480000 428.190000 ;
      RECT 0.000000 387.775000 1925.380000 388.675000 ;
      RECT 0.000000 381.380000 1926.480000 387.775000 ;
      RECT 1.100000 380.480000 1926.480000 381.380000 ;
      RECT 0.000000 340.100000 1926.480000 380.480000 ;
      RECT 0.000000 339.200000 1925.380000 340.100000 ;
      RECT 0.000000 333.760000 1926.480000 339.200000 ;
      RECT 1.100000 332.860000 1926.480000 333.760000 ;
      RECT 0.000000 291.715000 1926.480000 332.860000 ;
      RECT 0.000000 290.815000 1925.380000 291.715000 ;
      RECT 0.000000 286.050000 1926.480000 290.815000 ;
      RECT 1.100000 285.150000 1926.480000 286.050000 ;
      RECT 0.000000 242.945000 1926.480000 285.150000 ;
      RECT 0.000000 242.045000 1925.380000 242.945000 ;
      RECT 0.000000 238.435000 1926.480000 242.045000 ;
      RECT 1.100000 237.535000 1926.480000 238.435000 ;
      RECT 0.000000 194.465000 1926.480000 237.535000 ;
      RECT 0.000000 193.565000 1925.380000 194.465000 ;
      RECT 0.000000 190.720000 1926.480000 193.565000 ;
      RECT 1.100000 189.820000 1926.480000 190.720000 ;
      RECT 0.000000 145.985000 1926.480000 189.820000 ;
      RECT 0.000000 145.085000 1925.380000 145.985000 ;
      RECT 0.000000 143.105000 1926.480000 145.085000 ;
      RECT 1.100000 142.205000 1926.480000 143.105000 ;
      RECT 0.000000 97.315000 1926.480000 142.205000 ;
      RECT 0.000000 96.415000 1925.380000 97.315000 ;
      RECT 0.000000 95.490000 1926.480000 96.415000 ;
      RECT 1.100000 94.590000 1926.480000 95.490000 ;
      RECT 0.000000 48.545000 1926.480000 94.590000 ;
      RECT 0.000000 47.780000 1925.380000 48.545000 ;
      RECT 1.100000 47.645000 1925.380000 47.780000 ;
      RECT 1.100000 46.880000 1926.480000 47.645000 ;
      RECT 0.000000 17.460000 1926.480000 46.880000 ;
      RECT 1914.100000 12.660000 1926.480000 17.460000 ;
      RECT 0.000000 12.660000 12.380000 17.460000 ;
      RECT 0.000000 11.660000 1926.480000 12.660000 ;
      RECT 1919.900000 6.860000 1926.480000 11.660000 ;
      RECT 0.000000 6.860000 6.580000 11.660000 ;
      RECT 0.000000 2.465000 1926.480000 6.860000 ;
      RECT 0.000000 1.565000 1925.380000 2.465000 ;
      RECT 0.000000 1.220000 1926.480000 1.565000 ;
      RECT 1.100000 0.320000 1926.480000 1.220000 ;
      RECT 0.000000 0.000000 1926.480000 0.320000 ;
    LAYER met4 ;
      RECT 0.000000 2587.340000 1926.480000 2595.220000 ;
      RECT 11.380000 2581.540000 1915.100000 2587.340000 ;
      RECT 1914.100000 12.660000 1915.100000 2581.540000 ;
      RECT 17.180000 12.660000 1909.300000 2581.540000 ;
      RECT 11.380000 12.660000 12.380000 2581.540000 ;
      RECT 1919.900000 6.860000 1926.480000 2587.340000 ;
      RECT 11.380000 6.860000 1915.100000 12.660000 ;
      RECT 0.000000 6.860000 6.580000 2587.340000 ;
      RECT 0.000000 0.000000 1926.480000 6.860000 ;
  END
END rest_top

END LIBRARY
