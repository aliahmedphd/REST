##
## LEF for PtnCells ;
## created by Innovus v20.10-p004_1 on Mon Dec 27 16:42:06 2021
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO rest_top
  CLASS BLOCK ;
  SIZE 2369.460000 BY 2290.240000 ;
  FOREIGN rest_top 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1939 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 69.124 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 369.128 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.9548 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.248 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.982 LAYER met4  ;
    ANTENNAMAXAREACAR 55.4714 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 278.874 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.496244 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 4.530000 0.000000 4.670000 0.490000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.8133 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.8405 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 16.5434 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 81.5051 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1.930000 0.000000 2.070000 0.485000 ;
    END
  END wb_rst_i
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.530000 0.000000 496.670000 0.490000 ;
    END
  END wbs_stb_i
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.930000 0.000000 167.070000 0.490000 ;
    END
  END wbs_cyc_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.230000 0.000000 501.370000 0.490000 ;
    END
  END wbs_we_i
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.730000 0.000000 491.870000 0.490000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.930000 0.000000 487.070000 0.490000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.130000 0.000000 482.270000 0.490000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.430000 0.000000 477.570000 0.490000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.830000 0.000000 319.970000 0.490000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.030000 0.000000 315.170000 0.490000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.230000 0.000000 310.370000 0.490000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.430000 0.000000 305.570000 0.490000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.630000 0.000000 300.770000 0.490000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.830000 0.000000 295.970000 0.490000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.130000 0.000000 291.270000 0.490000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.430000 0.000000 286.570000 0.490000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.630000 0.000000 281.770000 0.490000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.830000 0.000000 276.970000 0.490000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.030000 0.000000 272.170000 0.490000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.230000 0.000000 267.370000 0.490000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.530000 0.000000 262.670000 0.490000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.730000 0.000000 257.870000 0.490000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.930000 0.000000 253.070000 0.490000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.130000 0.000000 248.270000 0.490000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.330000 0.000000 243.470000 0.490000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.630000 0.000000 238.770000 0.490000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.930000 0.000000 234.070000 0.490000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.030000 0.000000 229.170000 0.490000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.230000 0.000000 224.370000 0.490000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.430000 0.000000 219.570000 0.490000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.630000 0.000000 214.770000 0.490000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.830000 0.000000 209.970000 0.490000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.030000 0.000000 205.170000 0.490000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.330000 0.000000 200.470000 0.490000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.530000 0.000000 195.670000 0.490000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.830000 0.000000 190.970000 0.490000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.030000 0.000000 186.170000 0.490000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.230000 0.000000 181.370000 0.490000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.430000 0.000000 176.570000 0.490000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.730000 0.000000 171.870000 0.490000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.130000 0.000000 162.270000 0.490000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.330000 0.000000 157.470000 0.490000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.530000 0.000000 152.670000 0.490000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.730000 0.000000 147.870000 0.490000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.130000 0.000000 143.270000 0.490000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.330000 0.000000 138.470000 0.490000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.530000 0.000000 133.670000 0.490000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.730000 0.000000 128.870000 0.490000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.930000 0.000000 124.070000 0.490000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.130000 0.000000 119.270000 0.490000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.430000 0.000000 114.570000 0.490000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.630000 0.000000 109.770000 0.490000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.830000 0.000000 104.970000 0.490000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.030000 0.000000 100.170000 0.490000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.330000 0.000000 95.470000 0.490000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.530000 0.000000 90.670000 0.490000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.830000 0.000000 85.970000 0.490000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.030000 0.000000 81.170000 0.490000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.230000 0.000000 76.370000 0.490000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.430000 0.000000 71.570000 0.490000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.630000 0.000000 66.770000 0.490000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.830000 0.000000 61.970000 0.490000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130000 0.000000 57.270000 0.490000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.330000 0.000000 52.470000 0.490000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.630000 0.000000 47.770000 0.490000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.830000 0.000000 42.970000 0.490000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.030000 0.000000 38.170000 0.490000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.230000 0.000000 33.370000 0.490000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.530000 0.000000 28.670000 0.490000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.730000 0.000000 23.870000 0.490000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.930000 0.000000 19.070000 0.490000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.130000 0.000000 14.270000 0.490000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_ack_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9448 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.616 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 9.330000 0.000000 9.470000 0.490000 ;
    END
  END wbs_ack_o
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 472.630000 0.000000 472.770000 0.490000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 467.730000 0.000000 467.870000 0.490000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9252 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.518 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 463.030000 0.000000 463.170000 0.490000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.928 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.532 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 458.230000 0.000000 458.370000 0.490000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 453.430000 0.000000 453.570000 0.490000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8762 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.273 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 448.630000 0.000000 448.770000 0.490000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 443.830000 0.000000 443.970000 0.490000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9364 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.574 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 439.030000 0.000000 439.170000 0.490000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9707 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.7455 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 434.330000 0.000000 434.470000 0.490000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 429.630000 0.000000 429.770000 0.490000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 424.830000 0.000000 424.970000 0.490000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8874 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.329 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 420.030000 0.000000 420.170000 0.490000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9196 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.49 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 415.230000 0.000000 415.370000 0.490000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9336 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.56 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 410.430000 0.000000 410.570000 0.490000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9154 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.469 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 405.730000 0.000000 405.870000 0.490000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 400.930000 0.000000 401.070000 0.490000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 396.130000 0.000000 396.270000 0.490000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9126 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.455 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 391.330000 0.000000 391.470000 0.490000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9364 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.574 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 386.530000 0.000000 386.670000 0.490000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9182 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.483 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 381.830000 0.000000 381.970000 0.490000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 377.130000 0.000000 377.270000 0.490000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 372.330000 0.000000 372.470000 0.490000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 367.530000 0.000000 367.670000 0.490000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.928 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.532 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 362.730000 0.000000 362.870000 0.490000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9252 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.518 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 357.930000 0.000000 358.070000 0.490000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 353.130000 0.000000 353.270000 0.490000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 348.430000 0.000000 348.570000 0.490000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 343.630000 0.000000 343.770000 0.490000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8874 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.329 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 338.830000 0.000000 338.970000 0.490000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9392 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.588 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 334.130000 0.000000 334.270000 0.490000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 329.330000 0.000000 329.470000 0.490000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9266 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.525 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 324.530000 0.000000 324.670000 0.490000 ;
    END
  END wbs_dat_o[0]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1112.430000 0.000000 1112.570000 0.490000 ;
    END
  END la_data_in[127]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1107.730000 0.000000 1107.870000 0.490000 ;
    END
  END la_data_in[126]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1103.030000 0.000000 1103.170000 0.490000 ;
    END
  END la_data_in[125]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1098.230000 0.000000 1098.370000 0.490000 ;
    END
  END la_data_in[124]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1093.430000 0.000000 1093.570000 0.490000 ;
    END
  END la_data_in[123]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1088.630000 0.000000 1088.770000 0.490000 ;
    END
  END la_data_in[122]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1083.830000 0.000000 1083.970000 0.490000 ;
    END
  END la_data_in[121]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1079.130000 0.000000 1079.270000 0.490000 ;
    END
  END la_data_in[120]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1074.330000 0.000000 1074.470000 0.490000 ;
    END
  END la_data_in[119]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1069.530000 0.000000 1069.670000 0.490000 ;
    END
  END la_data_in[118]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1064.730000 0.000000 1064.870000 0.490000 ;
    END
  END la_data_in[117]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.930000 0.000000 1060.070000 0.490000 ;
    END
  END la_data_in[116]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1055.230000 0.000000 1055.370000 0.490000 ;
    END
  END la_data_in[115]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1050.530000 0.000000 1050.670000 0.490000 ;
    END
  END la_data_in[114]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1045.730000 0.000000 1045.870000 0.490000 ;
    END
  END la_data_in[113]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1040.930000 0.000000 1041.070000 0.490000 ;
    END
  END la_data_in[112]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.130000 0.000000 1036.270000 0.490000 ;
    END
  END la_data_in[111]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1031.330000 0.000000 1031.470000 0.490000 ;
    END
  END la_data_in[110]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1026.530000 0.000000 1026.670000 0.490000 ;
    END
  END la_data_in[109]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1021.830000 0.000000 1021.970000 0.490000 ;
    END
  END la_data_in[108]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1017.030000 0.000000 1017.170000 0.490000 ;
    END
  END la_data_in[107]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1012.230000 0.000000 1012.370000 0.490000 ;
    END
  END la_data_in[106]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.530000 0.000000 1007.670000 0.490000 ;
    END
  END la_data_in[105]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1002.730000 0.000000 1002.870000 0.490000 ;
    END
  END la_data_in[104]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 997.930000 0.000000 998.070000 0.490000 ;
    END
  END la_data_in[103]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 993.230000 0.000000 993.370000 0.490000 ;
    END
  END la_data_in[102]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 988.430000 0.000000 988.570000 0.490000 ;
    END
  END la_data_in[101]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 983.630000 0.000000 983.770000 0.490000 ;
    END
  END la_data_in[100]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.830000 0.000000 978.970000 0.490000 ;
    END
  END la_data_in[99]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 974.030000 0.000000 974.170000 0.490000 ;
    END
  END la_data_in[98]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 969.230000 0.000000 969.370000 0.490000 ;
    END
  END la_data_in[97]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 964.530000 0.000000 964.670000 0.490000 ;
    END
  END la_data_in[96]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.830000 0.000000 959.970000 0.490000 ;
    END
  END la_data_in[95]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 955.030000 0.000000 955.170000 0.490000 ;
    END
  END la_data_in[94]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 950.230000 0.000000 950.370000 0.490000 ;
    END
  END la_data_in[93]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 945.330000 0.000000 945.470000 0.490000 ;
    END
  END la_data_in[92]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 940.530000 0.000000 940.670000 0.490000 ;
    END
  END la_data_in[91]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 935.730000 0.000000 935.870000 0.490000 ;
    END
  END la_data_in[90]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 931.030000 0.000000 931.170000 0.490000 ;
    END
  END la_data_in[89]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 926.230000 0.000000 926.370000 0.490000 ;
    END
  END la_data_in[88]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.430000 0.000000 921.570000 0.490000 ;
    END
  END la_data_in[87]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 916.630000 0.000000 916.770000 0.490000 ;
    END
  END la_data_in[86]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.830000 0.000000 911.970000 0.490000 ;
    END
  END la_data_in[85]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.130000 0.000000 907.270000 0.490000 ;
    END
  END la_data_in[84]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 902.430000 0.000000 902.570000 0.490000 ;
    END
  END la_data_in[83]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 897.630000 0.000000 897.770000 0.490000 ;
    END
  END la_data_in[82]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.830000 0.000000 892.970000 0.490000 ;
    END
  END la_data_in[81]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.030000 0.000000 888.170000 0.490000 ;
    END
  END la_data_in[80]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 883.230000 0.000000 883.370000 0.490000 ;
    END
  END la_data_in[79]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 878.430000 0.000000 878.570000 0.490000 ;
    END
  END la_data_in[78]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 873.730000 0.000000 873.870000 0.490000 ;
    END
  END la_data_in[77]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 868.930000 0.000000 869.070000 0.490000 ;
    END
  END la_data_in[76]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 864.130000 0.000000 864.270000 0.490000 ;
    END
  END la_data_in[75]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.430000 0.000000 859.570000 0.490000 ;
    END
  END la_data_in[74]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 854.630000 0.000000 854.770000 0.490000 ;
    END
  END la_data_in[73]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 849.830000 0.000000 849.970000 0.490000 ;
    END
  END la_data_in[72]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 845.130000 0.000000 845.270000 0.490000 ;
    END
  END la_data_in[71]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.330000 0.000000 840.470000 0.490000 ;
    END
  END la_data_in[70]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.530000 0.000000 835.670000 0.490000 ;
    END
  END la_data_in[69]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.730000 0.000000 830.870000 0.490000 ;
    END
  END la_data_in[68]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 825.930000 0.000000 826.070000 0.490000 ;
    END
  END la_data_in[67]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.130000 0.000000 821.270000 0.490000 ;
    END
  END la_data_in[66]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 816.430000 0.000000 816.570000 0.490000 ;
    END
  END la_data_in[65]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.730000 0.000000 811.870000 0.490000 ;
    END
  END la_data_in[64]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.930000 0.000000 807.070000 0.490000 ;
    END
  END la_data_in[63]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 802.130000 0.000000 802.270000 0.490000 ;
    END
  END la_data_in[62]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.330000 0.000000 797.470000 0.490000 ;
    END
  END la_data_in[61]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.530000 0.000000 792.670000 0.490000 ;
    END
  END la_data_in[60]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 787.830000 0.000000 787.970000 0.490000 ;
    END
  END la_data_in[59]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.030000 0.000000 783.170000 0.490000 ;
    END
  END la_data_in[58]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 778.230000 0.000000 778.370000 0.490000 ;
    END
  END la_data_in[57]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 773.430000 0.000000 773.570000 0.490000 ;
    END
  END la_data_in[56]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 768.630000 0.000000 768.770000 0.490000 ;
    END
  END la_data_in[55]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.930000 0.000000 764.070000 0.490000 ;
    END
  END la_data_in[54]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 759.230000 0.000000 759.370000 0.490000 ;
    END
  END la_data_in[53]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.430000 0.000000 754.570000 0.490000 ;
    END
  END la_data_in[52]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.630000 0.000000 749.770000 0.490000 ;
    END
  END la_data_in[51]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 744.830000 0.000000 744.970000 0.490000 ;
    END
  END la_data_in[50]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.030000 0.000000 740.170000 0.490000 ;
    END
  END la_data_in[49]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.230000 0.000000 735.370000 0.490000 ;
    END
  END la_data_in[48]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.530000 0.000000 730.670000 0.490000 ;
    END
  END la_data_in[47]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.730000 0.000000 725.870000 0.490000 ;
    END
  END la_data_in[46]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.930000 0.000000 721.070000 0.490000 ;
    END
  END la_data_in[45]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.230000 0.000000 716.370000 0.490000 ;
    END
  END la_data_in[44]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.430000 0.000000 711.570000 0.490000 ;
    END
  END la_data_in[43]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.530000 0.000000 706.670000 0.490000 ;
    END
  END la_data_in[42]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 701.730000 0.000000 701.870000 0.490000 ;
    END
  END la_data_in[41]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.030000 0.000000 697.170000 0.490000 ;
    END
  END la_data_in[40]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.230000 0.000000 692.370000 0.490000 ;
    END
  END la_data_in[39]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 687.430000 0.000000 687.570000 0.490000 ;
    END
  END la_data_in[38]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.630000 0.000000 682.770000 0.490000 ;
    END
  END la_data_in[37]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 677.830000 0.000000 677.970000 0.490000 ;
    END
  END la_data_in[36]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.030000 0.000000 673.170000 0.490000 ;
    END
  END la_data_in[35]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.430000 0.000000 668.570000 0.490000 ;
    END
  END la_data_in[34]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.630000 0.000000 663.770000 0.490000 ;
    END
  END la_data_in[33]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.830000 0.000000 658.970000 0.490000 ;
    END
  END la_data_in[32]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 654.030000 0.000000 654.170000 0.490000 ;
    END
  END la_data_in[31]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.230000 0.000000 649.370000 0.490000 ;
    END
  END la_data_in[30]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.430000 0.000000 644.570000 0.490000 ;
    END
  END la_data_in[29]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.730000 0.000000 639.870000 0.490000 ;
    END
  END la_data_in[28]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.930000 0.000000 635.070000 0.490000 ;
    END
  END la_data_in[27]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.130000 0.000000 630.270000 0.490000 ;
    END
  END la_data_in[26]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 625.330000 0.000000 625.470000 0.490000 ;
    END
  END la_data_in[25]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.630000 0.000000 620.770000 0.490000 ;
    END
  END la_data_in[24]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.830000 0.000000 615.970000 0.490000 ;
    END
  END la_data_in[23]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.130000 0.000000 611.270000 0.490000 ;
    END
  END la_data_in[22]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.330000 0.000000 606.470000 0.490000 ;
    END
  END la_data_in[21]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601.530000 0.000000 601.670000 0.490000 ;
    END
  END la_data_in[20]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 596.730000 0.000000 596.870000 0.490000 ;
    END
  END la_data_in[19]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.930000 0.000000 592.070000 0.490000 ;
    END
  END la_data_in[18]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.130000 0.000000 587.270000 0.490000 ;
    END
  END la_data_in[17]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.430000 0.000000 582.570000 0.490000 ;
    END
  END la_data_in[16]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3956 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.87 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 30.1341 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 140.409 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 577.630000 0.000000 577.770000 0.490000 ;
    END
  END la_data_in[15]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.539 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 26.3234 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 121.909 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 572.930000 0.000000 573.070000 0.490000 ;
    END
  END la_data_in[14]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3956 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.87 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 32.3194 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 151.353 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 568.130000 0.000000 568.270000 0.490000 ;
    END
  END la_data_in[13]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0148 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.966 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 13.5465 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 65.7636 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 563.330000 0.000000 563.470000 0.490000 ;
    END
  END la_data_in[12]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4026 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.905 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 16.601 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 81.0364 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 558.530000 0.000000 558.670000 0.490000 ;
    END
  END la_data_in[11]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.0417 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.0475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.4348 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.456 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 49.9232 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 263.725 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 553.830000 0.000000 553.970000 0.490000 ;
    END
  END la_data_in[10]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9714 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.749 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 27.0528 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 125.02 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 549.030000 0.000000 549.170000 0.490000 ;
    END
  END la_data_in[9]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.5908 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.846 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 38.5495 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 189.655 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 544.230000 0.000000 544.370000 0.490000 ;
    END
  END la_data_in[8]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1222 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.503 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 18.3994 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 86.4505 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 539.430000 0.000000 539.570000 0.490000 ;
    END
  END la_data_in[7]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.355 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.667 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 14.5873 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 70.9677 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 534.630000 0.000000 534.770000 0.490000 ;
    END
  END la_data_in[6]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.1862 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.823 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 28.4331 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 138.531 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 529.830000 0.000000 529.970000 0.490000 ;
    END
  END la_data_in[5]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9928 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.738 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 21.8713 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 103.246 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 525.230000 0.000000 525.370000 0.490000 ;
    END
  END la_data_in[4]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9196 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.49 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 13.5893 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 63.0889 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 520.430000 0.000000 520.570000 0.490000 ;
    END
  END la_data_in[3]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0414 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.099 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 13.3202 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 64.6323 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 515.630000 0.000000 515.770000 0.490000 ;
    END
  END la_data_in[2]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5478 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.631 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 21.6279 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 102.624 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 510.830000 0.000000 510.970000 0.490000 ;
    END
  END la_data_in[1]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4138 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.961 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 16.7554 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 80.1111 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 506.030000 0.000000 506.170000 0.490000 ;
    END
  END la_data_in[0]
  PIN la_data_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9196 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.49 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1723.930000 0.000000 1724.070000 0.490000 ;
    END
  END la_data_out[127]
  PIN la_data_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9336 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.56 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1719.130000 0.000000 1719.270000 0.490000 ;
    END
  END la_data_out[126]
  PIN la_data_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1714.330000 0.000000 1714.470000 0.490000 ;
    END
  END la_data_out[125]
  PIN la_data_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1709.530000 0.000000 1709.670000 0.490000 ;
    END
  END la_data_out[124]
  PIN la_data_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1704.730000 0.000000 1704.870000 0.490000 ;
    END
  END la_data_out[123]
  PIN la_data_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9308 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.546 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1699.930000 0.000000 1700.070000 0.490000 ;
    END
  END la_data_out[122]
  PIN la_data_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9364 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.574 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1695.230000 0.000000 1695.370000 0.490000 ;
    END
  END la_data_out[121]
  PIN la_data_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.413 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1690.430000 0.000000 1690.570000 0.490000 ;
    END
  END la_data_out[120]
  PIN la_data_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1685.630000 0.000000 1685.770000 0.490000 ;
    END
  END la_data_out[119]
  PIN la_data_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1680.830000 0.000000 1680.970000 0.490000 ;
    END
  END la_data_out[118]
  PIN la_data_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9098 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.441 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1676.130000 0.000000 1676.270000 0.490000 ;
    END
  END la_data_out[117]
  PIN la_data_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1671.330000 0.000000 1671.470000 0.490000 ;
    END
  END la_data_out[116]
  PIN la_data_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1666.630000 0.000000 1666.770000 0.490000 ;
    END
  END la_data_out[115]
  PIN la_data_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.879 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.287 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1661.730000 0.000000 1661.870000 0.490000 ;
    END
  END la_data_out[114]
  PIN la_data_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1656.930000 0.000000 1657.070000 0.490000 ;
    END
  END la_data_out[113]
  PIN la_data_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9252 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.518 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1652.130000 0.000000 1652.270000 0.490000 ;
    END
  END la_data_out[112]
  PIN la_data_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.928 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.532 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1647.330000 0.000000 1647.470000 0.490000 ;
    END
  END la_data_out[111]
  PIN la_data_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1642.530000 0.000000 1642.670000 0.490000 ;
    END
  END la_data_out[110]
  PIN la_data_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1637.730000 0.000000 1637.870000 0.490000 ;
    END
  END la_data_out[109]
  PIN la_data_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8902 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1633.030000 0.000000 1633.170000 0.490000 ;
    END
  END la_data_out[108]
  PIN la_data_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1628.330000 0.000000 1628.470000 0.490000 ;
    END
  END la_data_out[107]
  PIN la_data_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1623.530000 0.000000 1623.670000 0.490000 ;
    END
  END la_data_out[106]
  PIN la_data_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1618.730000 0.000000 1618.870000 0.490000 ;
    END
  END la_data_out[105]
  PIN la_data_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1613.930000 0.000000 1614.070000 0.490000 ;
    END
  END la_data_out[104]
  PIN la_data_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1609.130000 0.000000 1609.270000 0.490000 ;
    END
  END la_data_out[103]
  PIN la_data_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1604.430000 0.000000 1604.570000 0.490000 ;
    END
  END la_data_out[102]
  PIN la_data_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1599.630000 0.000000 1599.770000 0.490000 ;
    END
  END la_data_out[101]
  PIN la_data_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1594.830000 0.000000 1594.970000 0.490000 ;
    END
  END la_data_out[100]
  PIN la_data_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1590.030000 0.000000 1590.170000 0.490000 ;
    END
  END la_data_out[99]
  PIN la_data_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.928 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.532 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1585.230000 0.000000 1585.370000 0.490000 ;
    END
  END la_data_out[98]
  PIN la_data_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1580.530000 0.000000 1580.670000 0.490000 ;
    END
  END la_data_out[97]
  PIN la_data_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1575.830000 0.000000 1575.970000 0.490000 ;
    END
  END la_data_out[96]
  PIN la_data_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1571.030000 0.000000 1571.170000 0.490000 ;
    END
  END la_data_out[95]
  PIN la_data_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.413 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1566.230000 0.000000 1566.370000 0.490000 ;
    END
  END la_data_out[94]
  PIN la_data_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1561.430000 0.000000 1561.570000 0.490000 ;
    END
  END la_data_out[93]
  PIN la_data_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1556.630000 0.000000 1556.770000 0.490000 ;
    END
  END la_data_out[92]
  PIN la_data_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.928 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.532 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1551.830000 0.000000 1551.970000 0.490000 ;
    END
  END la_data_out[91]
  PIN la_data_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1547.130000 0.000000 1547.270000 0.490000 ;
    END
  END la_data_out[90]
  PIN la_data_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.907 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.427 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1542.330000 0.000000 1542.470000 0.490000 ;
    END
  END la_data_out[89]
  PIN la_data_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.879 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.287 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1537.530000 0.000000 1537.670000 0.490000 ;
    END
  END la_data_out[88]
  PIN la_data_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9336 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.56 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1532.830000 0.000000 1532.970000 0.490000 ;
    END
  END la_data_out[87]
  PIN la_data_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1528.030000 0.000000 1528.170000 0.490000 ;
    END
  END la_data_out[86]
  PIN la_data_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9392 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.588 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1523.230000 0.000000 1523.370000 0.490000 ;
    END
  END la_data_out[85]
  PIN la_data_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1518.530000 0.000000 1518.670000 0.490000 ;
    END
  END la_data_out[84]
  PIN la_data_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1513.730000 0.000000 1513.870000 0.490000 ;
    END
  END la_data_out[83]
  PIN la_data_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9364 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.574 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1508.930000 0.000000 1509.070000 0.490000 ;
    END
  END la_data_out[82]
  PIN la_data_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1504.130000 0.000000 1504.270000 0.490000 ;
    END
  END la_data_out[81]
  PIN la_data_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1499.330000 0.000000 1499.470000 0.490000 ;
    END
  END la_data_out[80]
  PIN la_data_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1494.530000 0.000000 1494.670000 0.490000 ;
    END
  END la_data_out[79]
  PIN la_data_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1489.830000 0.000000 1489.970000 0.490000 ;
    END
  END la_data_out[78]
  PIN la_data_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.928 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.532 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1485.130000 0.000000 1485.270000 0.490000 ;
    END
  END la_data_out[77]
  PIN la_data_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9252 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.518 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1480.330000 0.000000 1480.470000 0.490000 ;
    END
  END la_data_out[76]
  PIN la_data_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1475.530000 0.000000 1475.670000 0.490000 ;
    END
  END la_data_out[75]
  PIN la_data_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1470.730000 0.000000 1470.870000 0.490000 ;
    END
  END la_data_out[74]
  PIN la_data_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1465.930000 0.000000 1466.070000 0.490000 ;
    END
  END la_data_out[73]
  PIN la_data_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9252 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.518 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1461.230000 0.000000 1461.370000 0.490000 ;
    END
  END la_data_out[72]
  PIN la_data_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.928 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.532 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1456.430000 0.000000 1456.570000 0.490000 ;
    END
  END la_data_out[71]
  PIN la_data_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1451.630000 0.000000 1451.770000 0.490000 ;
    END
  END la_data_out[70]
  PIN la_data_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1446.830000 0.000000 1446.970000 0.490000 ;
    END
  END la_data_out[69]
  PIN la_data_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.413 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1442.030000 0.000000 1442.170000 0.490000 ;
    END
  END la_data_out[68]
  PIN la_data_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9182 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.483 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1437.330000 0.000000 1437.470000 0.490000 ;
    END
  END la_data_out[67]
  PIN la_data_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9364 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.574 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1432.630000 0.000000 1432.770000 0.490000 ;
    END
  END la_data_out[66]
  PIN la_data_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8958 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.371 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1427.830000 0.000000 1427.970000 0.490000 ;
    END
  END la_data_out[65]
  PIN la_data_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1422.930000 0.000000 1423.070000 0.490000 ;
    END
  END la_data_out[64]
  PIN la_data_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1418.130000 0.000000 1418.270000 0.490000 ;
    END
  END la_data_out[63]
  PIN la_data_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.879 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.287 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1413.330000 0.000000 1413.470000 0.490000 ;
    END
  END la_data_out[62]
  PIN la_data_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9154 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.469 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1408.530000 0.000000 1408.670000 0.490000 ;
    END
  END la_data_out[61]
  PIN la_data_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1403.730000 0.000000 1403.870000 0.490000 ;
    END
  END la_data_out[60]
  PIN la_data_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9392 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.588 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1399.030000 0.000000 1399.170000 0.490000 ;
    END
  END la_data_out[59]
  PIN la_data_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1394.230000 0.000000 1394.370000 0.490000 ;
    END
  END la_data_out[58]
  PIN la_data_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1389.530000 0.000000 1389.670000 0.490000 ;
    END
  END la_data_out[57]
  PIN la_data_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9364 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.574 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1384.730000 0.000000 1384.870000 0.490000 ;
    END
  END la_data_out[56]
  PIN la_data_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1379.930000 0.000000 1380.070000 0.490000 ;
    END
  END la_data_out[55]
  PIN la_data_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1375.130000 0.000000 1375.270000 0.490000 ;
    END
  END la_data_out[54]
  PIN la_data_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1370.430000 0.000000 1370.570000 0.490000 ;
    END
  END la_data_out[53]
  PIN la_data_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1365.630000 0.000000 1365.770000 0.490000 ;
    END
  END la_data_out[52]
  PIN la_data_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9392 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.588 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1360.830000 0.000000 1360.970000 0.490000 ;
    END
  END la_data_out[51]
  PIN la_data_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1356.030000 0.000000 1356.170000 0.490000 ;
    END
  END la_data_out[50]
  PIN la_data_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1351.230000 0.000000 1351.370000 0.490000 ;
    END
  END la_data_out[49]
  PIN la_data_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1346.430000 0.000000 1346.570000 0.490000 ;
    END
  END la_data_out[48]
  PIN la_data_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1341.830000 0.000000 1341.970000 0.490000 ;
    END
  END la_data_out[47]
  PIN la_data_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9252 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.518 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1337.030000 0.000000 1337.170000 0.490000 ;
    END
  END la_data_out[46]
  PIN la_data_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.928 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.532 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1332.230000 0.000000 1332.370000 0.490000 ;
    END
  END la_data_out[45]
  PIN la_data_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1327.430000 0.000000 1327.570000 0.490000 ;
    END
  END la_data_out[44]
  PIN la_data_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1322.630000 0.000000 1322.770000 0.490000 ;
    END
  END la_data_out[43]
  PIN la_data_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.413 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1317.830000 0.000000 1317.970000 0.490000 ;
    END
  END la_data_out[42]
  PIN la_data_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9196 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.49 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1313.130000 0.000000 1313.270000 0.490000 ;
    END
  END la_data_out[41]
  PIN la_data_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1308.330000 0.000000 1308.470000 0.490000 ;
    END
  END la_data_out[40]
  PIN la_data_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8986 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.385 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1303.530000 0.000000 1303.670000 0.490000 ;
    END
  END la_data_out[39]
  PIN la_data_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1298.730000 0.000000 1298.870000 0.490000 ;
    END
  END la_data_out[38]
  PIN la_data_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1294.030000 0.000000 1294.170000 0.490000 ;
    END
  END la_data_out[37]
  PIN la_data_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.893 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.357 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1289.230000 0.000000 1289.370000 0.490000 ;
    END
  END la_data_out[36]
  PIN la_data_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1284.530000 0.000000 1284.670000 0.490000 ;
    END
  END la_data_out[35]
  PIN la_data_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1279.730000 0.000000 1279.870000 0.490000 ;
    END
  END la_data_out[34]
  PIN la_data_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9252 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.518 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1274.930000 0.000000 1275.070000 0.490000 ;
    END
  END la_data_out[33]
  PIN la_data_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1270.130000 0.000000 1270.270000 0.490000 ;
    END
  END la_data_out[32]
  PIN la_data_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1265.330000 0.000000 1265.470000 0.490000 ;
    END
  END la_data_out[31]
  PIN la_data_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1260.530000 0.000000 1260.670000 0.490000 ;
    END
  END la_data_out[30]
  PIN la_data_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1255.830000 0.000000 1255.970000 0.490000 ;
    END
  END la_data_out[29]
  PIN la_data_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1251.030000 0.000000 1251.170000 0.490000 ;
    END
  END la_data_out[28]
  PIN la_data_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9364 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.574 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1246.330000 0.000000 1246.470000 0.490000 ;
    END
  END la_data_out[27]
  PIN la_data_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1241.530000 0.000000 1241.670000 0.490000 ;
    END
  END la_data_out[26]
  PIN la_data_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1236.730000 0.000000 1236.870000 0.490000 ;
    END
  END la_data_out[25]
  PIN la_data_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1231.930000 0.000000 1232.070000 0.490000 ;
    END
  END la_data_out[24]
  PIN la_data_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1227.230000 0.000000 1227.370000 0.490000 ;
    END
  END la_data_out[23]
  PIN la_data_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9336 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.56 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1222.430000 0.000000 1222.570000 0.490000 ;
    END
  END la_data_out[22]
  PIN la_data_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9154 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.469 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1217.630000 0.000000 1217.770000 0.490000 ;
    END
  END la_data_out[21]
  PIN la_data_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1212.830000 0.000000 1212.970000 0.490000 ;
    END
  END la_data_out[20]
  PIN la_data_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8846 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.315 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1208.030000 0.000000 1208.170000 0.490000 ;
    END
  END la_data_out[19]
  PIN la_data_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1203.230000 0.000000 1203.370000 0.490000 ;
    END
  END la_data_out[18]
  PIN la_data_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1198.630000 0.000000 1198.770000 0.490000 ;
    END
  END la_data_out[17]
  PIN la_data_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9364 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.574 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1193.830000 0.000000 1193.970000 0.490000 ;
    END
  END la_data_out[16]
  PIN la_data_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1189.030000 0.000000 1189.170000 0.490000 ;
    END
  END la_data_out[15]
  PIN la_data_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1184.130000 0.000000 1184.270000 0.490000 ;
    END
  END la_data_out[14]
  PIN la_data_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8986 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.385 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1179.330000 0.000000 1179.470000 0.490000 ;
    END
  END la_data_out[13]
  PIN la_data_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9392 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.588 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1174.530000 0.000000 1174.670000 0.490000 ;
    END
  END la_data_out[12]
  PIN la_data_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1169.730000 0.000000 1169.870000 0.490000 ;
    END
  END la_data_out[11]
  PIN la_data_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.893 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.357 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1165.030000 0.000000 1165.170000 0.490000 ;
    END
  END la_data_out[10]
  PIN la_data_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1160.230000 0.000000 1160.370000 0.490000 ;
    END
  END la_data_out[9]
  PIN la_data_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1155.430000 0.000000 1155.570000 0.490000 ;
    END
  END la_data_out[8]
  PIN la_data_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9252 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.518 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1150.730000 0.000000 1150.870000 0.490000 ;
    END
  END la_data_out[7]
  PIN la_data_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.928 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.532 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1145.930000 0.000000 1146.070000 0.490000 ;
    END
  END la_data_out[6]
  PIN la_data_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1141.130000 0.000000 1141.270000 0.490000 ;
    END
  END la_data_out[5]
  PIN la_data_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1136.430000 0.000000 1136.570000 0.490000 ;
    END
  END la_data_out[4]
  PIN la_data_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1131.630000 0.000000 1131.770000 0.490000 ;
    END
  END la_data_out[3]
  PIN la_data_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9182 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.483 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1126.830000 0.000000 1126.970000 0.490000 ;
    END
  END la_data_out[2]
  PIN la_data_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9308 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.546 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1122.030000 0.000000 1122.170000 0.490000 ;
    END
  END la_data_out[1]
  PIN la_data_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1117.230000 0.000000 1117.370000 0.490000 ;
    END
  END la_data_out[0]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2335.130000 0.000000 2335.270000 0.490000 ;
    END
  END la_oenb[127]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2330.330000 0.000000 2330.470000 0.490000 ;
    END
  END la_oenb[126]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2325.530000 0.000000 2325.670000 0.490000 ;
    END
  END la_oenb[125]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2320.730000 0.000000 2320.870000 0.490000 ;
    END
  END la_oenb[124]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2315.930000 0.000000 2316.070000 0.490000 ;
    END
  END la_oenb[123]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2311.130000 0.000000 2311.270000 0.490000 ;
    END
  END la_oenb[122]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2306.430000 0.000000 2306.570000 0.490000 ;
    END
  END la_oenb[121]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2301.730000 0.000000 2301.870000 0.490000 ;
    END
  END la_oenb[120]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2296.930000 0.000000 2297.070000 0.490000 ;
    END
  END la_oenb[119]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2292.130000 0.000000 2292.270000 0.490000 ;
    END
  END la_oenb[118]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2287.330000 0.000000 2287.470000 0.490000 ;
    END
  END la_oenb[117]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2282.530000 0.000000 2282.670000 0.490000 ;
    END
  END la_oenb[116]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2277.830000 0.000000 2277.970000 0.490000 ;
    END
  END la_oenb[115]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2273.030000 0.000000 2273.170000 0.490000 ;
    END
  END la_oenb[114]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2268.230000 0.000000 2268.370000 0.490000 ;
    END
  END la_oenb[113]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2263.430000 0.000000 2263.570000 0.490000 ;
    END
  END la_oenb[112]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2258.630000 0.000000 2258.770000 0.490000 ;
    END
  END la_oenb[111]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2253.930000 0.000000 2254.070000 0.490000 ;
    END
  END la_oenb[110]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2249.230000 0.000000 2249.370000 0.490000 ;
    END
  END la_oenb[109]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2244.430000 0.000000 2244.570000 0.490000 ;
    END
  END la_oenb[108]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2239.630000 0.000000 2239.770000 0.490000 ;
    END
  END la_oenb[107]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2234.830000 0.000000 2234.970000 0.490000 ;
    END
  END la_oenb[106]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2230.030000 0.000000 2230.170000 0.490000 ;
    END
  END la_oenb[105]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2225.230000 0.000000 2225.370000 0.490000 ;
    END
  END la_oenb[104]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2220.530000 0.000000 2220.670000 0.490000 ;
    END
  END la_oenb[103]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2215.730000 0.000000 2215.870000 0.490000 ;
    END
  END la_oenb[102]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2210.930000 0.000000 2211.070000 0.490000 ;
    END
  END la_oenb[101]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2206.230000 0.000000 2206.370000 0.490000 ;
    END
  END la_oenb[100]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2201.430000 0.000000 2201.570000 0.490000 ;
    END
  END la_oenb[99]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2196.630000 0.000000 2196.770000 0.490000 ;
    END
  END la_oenb[98]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2191.930000 0.000000 2192.070000 0.490000 ;
    END
  END la_oenb[97]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2187.130000 0.000000 2187.270000 0.490000 ;
    END
  END la_oenb[96]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2182.330000 0.000000 2182.470000 0.490000 ;
    END
  END la_oenb[95]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2177.530000 0.000000 2177.670000 0.490000 ;
    END
  END la_oenb[94]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2172.730000 0.000000 2172.870000 0.490000 ;
    END
  END la_oenb[93]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2167.930000 0.000000 2168.070000 0.490000 ;
    END
  END la_oenb[92]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2163.230000 0.000000 2163.370000 0.490000 ;
    END
  END la_oenb[91]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2158.530000 0.000000 2158.670000 0.490000 ;
    END
  END la_oenb[90]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2153.730000 0.000000 2153.870000 0.490000 ;
    END
  END la_oenb[89]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2148.930000 0.000000 2149.070000 0.490000 ;
    END
  END la_oenb[88]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2144.130000 0.000000 2144.270000 0.490000 ;
    END
  END la_oenb[87]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2139.230000 0.000000 2139.370000 0.490000 ;
    END
  END la_oenb[86]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2134.530000 0.000000 2134.670000 0.490000 ;
    END
  END la_oenb[85]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2129.730000 0.000000 2129.870000 0.490000 ;
    END
  END la_oenb[84]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2124.930000 0.000000 2125.070000 0.490000 ;
    END
  END la_oenb[83]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2120.130000 0.000000 2120.270000 0.490000 ;
    END
  END la_oenb[82]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2115.330000 0.000000 2115.470000 0.490000 ;
    END
  END la_oenb[81]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2110.530000 0.000000 2110.670000 0.490000 ;
    END
  END la_oenb[80]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2105.930000 0.000000 2106.070000 0.490000 ;
    END
  END la_oenb[79]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2101.130000 0.000000 2101.270000 0.490000 ;
    END
  END la_oenb[78]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2096.330000 0.000000 2096.470000 0.490000 ;
    END
  END la_oenb[77]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2091.530000 0.000000 2091.670000 0.490000 ;
    END
  END la_oenb[76]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2086.730000 0.000000 2086.870000 0.490000 ;
    END
  END la_oenb[75]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2081.930000 0.000000 2082.070000 0.490000 ;
    END
  END la_oenb[74]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2077.130000 0.000000 2077.270000 0.490000 ;
    END
  END la_oenb[73]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2072.430000 0.000000 2072.570000 0.490000 ;
    END
  END la_oenb[72]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2067.630000 0.000000 2067.770000 0.490000 ;
    END
  END la_oenb[71]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2062.830000 0.000000 2062.970000 0.490000 ;
    END
  END la_oenb[70]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2058.130000 0.000000 2058.270000 0.490000 ;
    END
  END la_oenb[69]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2053.330000 0.000000 2053.470000 0.490000 ;
    END
  END la_oenb[68]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2048.530000 0.000000 2048.670000 0.490000 ;
    END
  END la_oenb[67]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2043.830000 0.000000 2043.970000 0.490000 ;
    END
  END la_oenb[66]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2039.030000 0.000000 2039.170000 0.490000 ;
    END
  END la_oenb[65]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2034.230000 0.000000 2034.370000 0.490000 ;
    END
  END la_oenb[64]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2029.430000 0.000000 2029.570000 0.490000 ;
    END
  END la_oenb[63]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2024.630000 0.000000 2024.770000 0.490000 ;
    END
  END la_oenb[62]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2019.830000 0.000000 2019.970000 0.490000 ;
    END
  END la_oenb[61]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2015.130000 0.000000 2015.270000 0.490000 ;
    END
  END la_oenb[60]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2010.430000 0.000000 2010.570000 0.490000 ;
    END
  END la_oenb[59]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2005.630000 0.000000 2005.770000 0.490000 ;
    END
  END la_oenb[58]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2000.830000 0.000000 2000.970000 0.490000 ;
    END
  END la_oenb[57]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1996.030000 0.000000 1996.170000 0.490000 ;
    END
  END la_oenb[56]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1991.230000 0.000000 1991.370000 0.490000 ;
    END
  END la_oenb[55]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1986.530000 0.000000 1986.670000 0.490000 ;
    END
  END la_oenb[54]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1981.730000 0.000000 1981.870000 0.490000 ;
    END
  END la_oenb[53]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1976.930000 0.000000 1977.070000 0.490000 ;
    END
  END la_oenb[52]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1972.130000 0.000000 1972.270000 0.490000 ;
    END
  END la_oenb[51]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1967.330000 0.000000 1967.470000 0.490000 ;
    END
  END la_oenb[50]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1962.630000 0.000000 1962.770000 0.490000 ;
    END
  END la_oenb[49]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1957.930000 0.000000 1958.070000 0.490000 ;
    END
  END la_oenb[48]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1953.130000 0.000000 1953.270000 0.490000 ;
    END
  END la_oenb[47]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1948.330000 0.000000 1948.470000 0.490000 ;
    END
  END la_oenb[46]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1943.530000 0.000000 1943.670000 0.490000 ;
    END
  END la_oenb[45]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1938.730000 0.000000 1938.870000 0.490000 ;
    END
  END la_oenb[44]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1933.930000 0.000000 1934.070000 0.490000 ;
    END
  END la_oenb[43]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1929.230000 0.000000 1929.370000 0.490000 ;
    END
  END la_oenb[42]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1924.430000 0.000000 1924.570000 0.490000 ;
    END
  END la_oenb[41]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1919.630000 0.000000 1919.770000 0.490000 ;
    END
  END la_oenb[40]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1914.930000 0.000000 1915.070000 0.490000 ;
    END
  END la_oenb[39]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1910.130000 0.000000 1910.270000 0.490000 ;
    END
  END la_oenb[38]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.330000 0.000000 1905.470000 0.490000 ;
    END
  END la_oenb[37]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1900.530000 0.000000 1900.670000 0.490000 ;
    END
  END la_oenb[36]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1895.730000 0.000000 1895.870000 0.490000 ;
    END
  END la_oenb[35]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1890.930000 0.000000 1891.070000 0.490000 ;
    END
  END la_oenb[34]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1886.130000 0.000000 1886.270000 0.490000 ;
    END
  END la_oenb[33]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1881.330000 0.000000 1881.470000 0.490000 ;
    END
  END la_oenb[32]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1876.530000 0.000000 1876.670000 0.490000 ;
    END
  END la_oenb[31]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1871.730000 0.000000 1871.870000 0.490000 ;
    END
  END la_oenb[30]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1867.130000 0.000000 1867.270000 0.490000 ;
    END
  END la_oenb[29]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1862.330000 0.000000 1862.470000 0.490000 ;
    END
  END la_oenb[28]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1857.530000 0.000000 1857.670000 0.490000 ;
    END
  END la_oenb[27]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1852.730000 0.000000 1852.870000 0.490000 ;
    END
  END la_oenb[26]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1847.930000 0.000000 1848.070000 0.490000 ;
    END
  END la_oenb[25]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1843.130000 0.000000 1843.270000 0.490000 ;
    END
  END la_oenb[24]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1838.430000 0.000000 1838.570000 0.490000 ;
    END
  END la_oenb[23]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1833.630000 0.000000 1833.770000 0.490000 ;
    END
  END la_oenb[22]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1828.830000 0.000000 1828.970000 0.490000 ;
    END
  END la_oenb[21]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1824.030000 0.000000 1824.170000 0.490000 ;
    END
  END la_oenb[20]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1819.330000 0.000000 1819.470000 0.490000 ;
    END
  END la_oenb[19]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1814.530000 0.000000 1814.670000 0.490000 ;
    END
  END la_oenb[18]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1809.830000 0.000000 1809.970000 0.490000 ;
    END
  END la_oenb[17]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1805.030000 0.000000 1805.170000 0.490000 ;
    END
  END la_oenb[16]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1800.230000 0.000000 1800.370000 0.490000 ;
    END
  END la_oenb[15]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1795.430000 0.000000 1795.570000 0.490000 ;
    END
  END la_oenb[14]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1790.630000 0.000000 1790.770000 0.490000 ;
    END
  END la_oenb[13]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1785.830000 0.000000 1785.970000 0.490000 ;
    END
  END la_oenb[12]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1781.130000 0.000000 1781.270000 0.490000 ;
    END
  END la_oenb[11]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1776.330000 0.000000 1776.470000 0.490000 ;
    END
  END la_oenb[10]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1771.630000 0.000000 1771.770000 0.490000 ;
    END
  END la_oenb[9]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1766.830000 0.000000 1766.970000 0.490000 ;
    END
  END la_oenb[8]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1762.030000 0.000000 1762.170000 0.490000 ;
    END
  END la_oenb[7]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1757.230000 0.000000 1757.370000 0.490000 ;
    END
  END la_oenb[6]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1752.530000 0.000000 1752.670000 0.490000 ;
    END
  END la_oenb[5]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1747.730000 0.000000 1747.870000 0.490000 ;
    END
  END la_oenb[4]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1742.930000 0.000000 1743.070000 0.490000 ;
    END
  END la_oenb[3]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1738.130000 0.000000 1738.270000 0.490000 ;
    END
  END la_oenb[2]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1733.330000 0.000000 1733.470000 0.490000 ;
    END
  END la_oenb[1]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1728.530000 0.000000 1728.670000 0.490000 ;
    END
  END la_oenb[0]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 83.735000 0.800000 84.035000 ;
    END
  END io_in[37]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.1448 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.576 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 43.8601 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 214.862 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 2.6214 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.424 LAYER met3  ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 9.63176 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 31.566 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 209.800000 0.800000 210.100000 ;
    END
  END io_in[36]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4809 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.56 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.318 LAYER met3  ;
    ANTENNAMAXAREACAR 31.3148 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 153.978 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.287421 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 335.865000 0.800000 336.165000 ;
    END
  END io_in[35]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 504.300000 0.800000 504.600000 ;
    END
  END io_in[34]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 48.7819 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 260.632 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.1735 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 149.312 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 796.8 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.37 LAYER met4  ;
    ANTENNAMAXAREACAR 68.5579 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 349.012 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.409837 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 672.355000 0.800000 672.655000 ;
    END
  END io_in[33]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 41.0734 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 219.52 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.1735 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 150.02 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 801.52 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.2995 LAYER met4  ;
    ANTENNAMAXAREACAR 70.3389 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 356.901 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.286759 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 840.600000 0.800000 840.900000 ;
    END
  END io_in[32]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8759 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.448 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.1578 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 33.312 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 20.5509 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 103.635 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.460202 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1008.845000 0.800000 1009.145000 ;
    END
  END io_in[31]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.1578 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 33.312 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met4  ;
    ANTENNAMAXAREACAR 11.6495 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 59.1252 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.500049 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1176.900000 0.800000 1177.200000 ;
    END
  END io_in[30]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0629 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.144 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 5.36754 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 26.5845 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1345.145000 0.800000 1345.445000 ;
    END
  END io_in[29]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0948 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.304 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.9618 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 21.6 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 37.4244 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 195.394 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1513.485000 0.800000 1513.785000 ;
    END
  END io_in[28]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5964 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.656 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 5.27663 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 25.7791 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1681.540000 0.800000 1681.840000 ;
    END
  END io_in[27]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5904 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.624 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 5.30572 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 25.7643 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1849.880000 0.800000 1850.180000 ;
    END
  END io_in[26]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.6082 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3024 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.088 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8212 LAYER met3  ;
    ANTENNAMAXAREACAR 86.095 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 412.505 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.172915 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2018.030000 0.800000 2018.330000 ;
    END
  END io_in[25]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1574 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.616 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.1448 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.576 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 21.3149 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 111.507 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2186.180000 0.800000 2186.480000 ;
    END
  END io_in[24]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.330000 2289.750000 134.470000 2290.240000 ;
    END
  END io_in[23]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.530000 2289.750000 403.670000 2290.240000 ;
    END
  END io_in[22]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.530000 2289.750000 672.670000 2290.240000 ;
    END
  END io_in[21]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 941.730000 2289.750000 941.870000 2290.240000 ;
    END
  END io_in[20]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1210.830000 2289.750000 1210.970000 2290.240000 ;
    END
  END io_in[19]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1480.030000 2289.750000 1480.170000 2290.240000 ;
    END
  END io_in[18]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1749.130000 2289.750000 1749.270000 2290.240000 ;
    END
  END io_in[17]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2018.330000 2289.750000 2018.470000 2290.240000 ;
    END
  END io_in[16]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2287.430000 2289.750000 2287.570000 2290.240000 ;
    END
  END io_in[15]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 2142.575000 2369.460000 2142.875000 ;
    END
  END io_in[14]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 1971.005000 2369.460000 1971.305000 ;
    END
  END io_in[13]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 1799.625000 2369.460000 1799.925000 ;
    END
  END io_in[12]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 1628.245000 2369.460000 1628.545000 ;
    END
  END io_in[11]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 1456.675000 2369.460000 1456.975000 ;
    END
  END io_in[10]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 1285.390000 2369.460000 1285.690000 ;
    END
  END io_in[9]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.1448 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.576 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9555 LAYER met4  ;
    ANTENNAMAXAREACAR 16.4458 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 82.1642 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.382312 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 5.5089 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.824 LAYER met3  ;
    ANTENNAGATEAREA 0.9555 LAYER met3  ;
    ANTENNAMAXAREACAR 79.2681 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 386.635 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.283177 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 1113.915000 2369.460000 1114.215000 ;
    END
  END io_in[8]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 942.440000 2369.460000 942.740000 ;
    END
  END io_in[7]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 770.965000 2369.460000 771.265000 ;
    END
  END io_in[6]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6433 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.896 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.1448 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.576 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 33.1883 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 173.323 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 642.430000 2369.460000 642.730000 ;
    END
  END io_in[5]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 513.895000 2369.460000 514.195000 ;
    END
  END io_in[4]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 385.360000 2369.460000 385.660000 ;
    END
  END io_in[3]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 256.730000 2369.460000 257.030000 ;
    END
  END io_in[2]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 128.100000 2369.460000 128.400000 ;
    END
  END io_in[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 2.415000 2369.460000 2.715000 ;
    END
  END io_in[0]
  PIN io_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.672 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 41.650000 0.800000 41.950000 ;
    END
  END io_out[37]
  PIN io_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2019 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.072 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 167.715000 0.800000 168.015000 ;
    END
  END io_out[36]
  PIN io_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0964 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.176 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 293.970000 0.800000 294.270000 ;
    END
  END io_out[35]
  PIN io_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.6544 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.152 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 462.120000 0.800000 462.420000 ;
    END
  END io_out[34]
  PIN io_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.3044 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 38.952 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 630.270000 0.800000 630.570000 ;
    END
  END io_out[33]
  PIN io_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.8669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.952 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 798.515000 0.800000 798.815000 ;
    END
  END io_out[32]
  PIN io_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.3144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.672 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 966.760000 0.800000 967.060000 ;
    END
  END io_out[31]
  PIN io_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.7304 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.024 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 63.0708 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 336.848 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1134.910000 0.800000 1135.210000 ;
    END
  END io_out[30]
  PIN io_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 152.741 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 815.088 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.3749 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.128 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1303.155000 0.800000 1303.455000 ;
    END
  END io_out[29]
  PIN io_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3579 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.904 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1471.305000 0.800000 1471.605000 ;
    END
  END io_out[28]
  PIN io_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.7905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 53.152 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1639.455000 0.800000 1639.755000 ;
    END
  END io_out[27]
  PIN io_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.5679 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.824 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.0858 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 48.928 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1807.795000 0.800000 1808.095000 ;
    END
  END io_out[26]
  PIN io_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6234 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.32 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1976.040000 0.800000 1976.340000 ;
    END
  END io_out[25]
  PIN io_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3314 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.096 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2144.190000 0.800000 2144.490000 ;
    END
  END io_out[24]
  PIN io_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.03 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 67.030000 2289.750000 67.170000 2290.240000 ;
    END
  END io_out[23]
  PIN io_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4696 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.122 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 336.230000 2289.750000 336.370000 2290.240000 ;
    END
  END io_out[22]
  PIN io_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 605.330000 2289.750000 605.470000 2290.240000 ;
    END
  END io_out[21]
  PIN io_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2302 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.925 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 874.430000 2289.750000 874.570000 2290.240000 ;
    END
  END io_out[20]
  PIN io_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1574 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.679 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1143.530000 2289.750000 1143.670000 2290.240000 ;
    END
  END io_out[19]
  PIN io_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.234 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.944 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1412.730000 2289.750000 1412.870000 2290.240000 ;
    END
  END io_out[18]
  PIN io_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.24 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.092 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1681.830000 2289.750000 1681.970000 2290.240000 ;
    END
  END io_out[17]
  PIN io_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.107 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.427 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1950.930000 2289.750000 1951.070000 2290.240000 ;
    END
  END io_out[16]
  PIN io_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.275 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.149 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2220.030000 2289.750000 2220.170000 2290.240000 ;
    END
  END io_out[15]
  PIN io_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5784 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.08 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 2185.420000 2369.460000 2185.720000 ;
    END
  END io_out[14]
  PIN io_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.0389 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.536 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 2013.945000 2369.460000 2014.245000 ;
    END
  END io_out[13]
  PIN io_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.5947 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 46.304 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 1842.565000 2369.460000 1842.865000 ;
    END
  END io_out[12]
  PIN io_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0674 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.688 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 1671.090000 2369.460000 1671.390000 ;
    END
  END io_out[11]
  PIN io_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.4909 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.08 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 13.5018 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 72.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 1499.615000 2369.460000 1499.915000 ;
    END
  END io_out[10]
  PIN io_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3024 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.608 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 1328.330000 2369.460000 1328.630000 ;
    END
  END io_out[9]
  PIN io_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.5789 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 46.216 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 66.9378 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 357.472 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 1156.855000 2369.460000 1157.155000 ;
    END
  END io_out[8]
  PIN io_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.496 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 985.380000 2369.460000 985.680000 ;
    END
  END io_out[7]
  PIN io_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.0774 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.888 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 814.000000 2369.460000 814.300000 ;
    END
  END io_out[6]
  PIN io_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.9844 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.912 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 685.370000 2369.460000 685.670000 ;
    END
  END io_out[5]
  PIN io_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.3939 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.096 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 556.645000 2369.460000 556.945000 ;
    END
  END io_out[4]
  PIN io_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.1329 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.704 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 428.205000 2369.460000 428.505000 ;
    END
  END io_out[3]
  PIN io_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2319 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.232 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 299.575000 2369.460000 299.875000 ;
    END
  END io_out[2]
  PIN io_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3219 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.712 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 170.945000 2369.460000 171.245000 ;
    END
  END io_out[1]
  PIN io_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2409 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.28 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 42.505000 2369.460000 42.805000 ;
    END
  END io_out[0]
  PIN io_oeb[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3849 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.048 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1.655000 0.800000 1.955000 ;
    END
  END io_oeb[37]
  PIN io_oeb[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3054 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.104 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 125.820000 0.800000 126.120000 ;
    END
  END io_oeb[36]
  PIN io_oeb[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2844 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.992 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 251.980000 0.800000 252.280000 ;
    END
  END io_oeb[35]
  PIN io_oeb[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2304 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.224 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 420.130000 0.800000 420.430000 ;
    END
  END io_oeb[34]
  PIN io_oeb[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.2582 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 55.176 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 588.280000 0.800000 588.580000 ;
    END
  END io_oeb[33]
  PIN io_oeb[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9234 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.92 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 756.430000 0.800000 756.730000 ;
    END
  END io_oeb[32]
  PIN io_oeb[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.2819 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 38.832 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 924.675000 0.800000 924.975000 ;
    END
  END io_oeb[31]
  PIN io_oeb[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8334 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.44 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1092.920000 0.800000 1093.220000 ;
    END
  END io_oeb[30]
  PIN io_oeb[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4664 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.816 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1261.070000 0.800000 1261.370000 ;
    END
  END io_oeb[29]
  PIN io_oeb[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1514 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.136 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1429.410000 0.800000 1429.710000 ;
    END
  END io_oeb[28]
  PIN io_oeb[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 33.9738 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 181.664 LAYER met4  ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.8509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1597.465000 0.800000 1597.765000 ;
    END
  END io_oeb[27]
  PIN io_oeb[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.7524 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.008 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1765.710000 0.800000 1766.010000 ;
    END
  END io_oeb[26]
  PIN io_oeb[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.2064 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.096 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1933.860000 0.800000 1934.160000 ;
    END
  END io_oeb[25]
  PIN io_oeb[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3969 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.592 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2102.105000 0.800000 2102.405000 ;
    END
  END io_oeb[24]
  PIN io_oeb[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1154 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.469 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 4.730000 2289.755000 4.870000 2290.240000 ;
    END
  END io_oeb[23]
  PIN io_oeb[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.8098 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.823 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 268.930000 2289.750000 269.070000 2290.240000 ;
    END
  END io_oeb[22]
  PIN io_oeb[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0946 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.365 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 538.130000 2289.750000 538.270000 2290.240000 ;
    END
  END io_oeb[21]
  PIN io_oeb[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8264 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.906 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 807.230000 2289.750000 807.370000 2290.240000 ;
    END
  END io_oeb[20]
  PIN io_oeb[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5648 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.598 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1076.330000 2289.750000 1076.470000 2290.240000 ;
    END
  END io_oeb[19]
  PIN io_oeb[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1518 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.651 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1345.430000 2289.750000 1345.570000 2290.240000 ;
    END
  END io_oeb[18]
  PIN io_oeb[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3058 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.303 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1614.630000 2289.750000 1614.770000 2290.240000 ;
    END
  END io_oeb[17]
  PIN io_oeb[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9658 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.721 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1883.730000 2289.750000 1883.870000 2290.240000 ;
    END
  END io_oeb[16]
  PIN io_oeb[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.184 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.694 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2152.830000 2289.750000 2152.970000 2290.240000 ;
    END
  END io_oeb[15]
  PIN io_oeb[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1769 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.272 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 2225.225000 2369.460000 2225.525000 ;
    END
  END io_oeb[14]
  PIN io_oeb[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9849 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.248 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 2056.885000 2369.460000 2057.185000 ;
    END
  END io_oeb[13]
  PIN io_oeb[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 21.2419 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 113.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 14.0268 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 75.28 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 1885.315000 2369.460000 1885.615000 ;
    END
  END io_oeb[12]
  PIN io_oeb[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8389 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 68.4018 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 365.28 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 1713.935000 2369.460000 1714.235000 ;
    END
  END io_oeb[11]
  PIN io_oeb[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.9374 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.128 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 45.8688 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 245.104 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 1542.460000 2369.460000 1542.760000 ;
    END
  END io_oeb[10]
  PIN io_oeb[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2424 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.288 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 1371.080000 2369.460000 1371.380000 ;
    END
  END io_oeb[9]
  PIN io_oeb[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5994 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.192 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 1199.700000 2369.460000 1200.000000 ;
    END
  END io_oeb[8]
  PIN io_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.4632 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.936 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 1028.320000 2369.460000 1028.620000 ;
    END
  END io_oeb[7]
  PIN io_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.6939 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.696 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 856.845000 2369.460000 857.145000 ;
    END
  END io_oeb[6]
  PIN io_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7839 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.176 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 728.215000 2369.460000 728.515000 ;
    END
  END io_oeb[5]
  PIN io_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.3169 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.352 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 599.585000 2369.460000 599.885000 ;
    END
  END io_oeb[4]
  PIN io_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2514 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.336 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 471.050000 2369.460000 471.350000 ;
    END
  END io_oeb[3]
  PIN io_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3039 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.616 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 342.515000 2369.460000 342.815000 ;
    END
  END io_oeb[2]
  PIN io_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2499 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 213.885000 2369.460000 214.185000 ;
    END
  END io_oeb[1]
  PIN io_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2259 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 85.255000 2369.460000 85.555000 ;
    END
  END io_oeb[0]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 378.045000 0.800000 378.345000 ;
    END
  END analog_io[28]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 546.290000 0.800000 546.590000 ;
    END
  END analog_io[27]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 714.535000 0.800000 714.835000 ;
    END
  END analog_io[26]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 882.590000 0.800000 882.890000 ;
    END
  END analog_io[25]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1050.835000 0.800000 1051.135000 ;
    END
  END analog_io[24]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1219.080000 0.800000 1219.380000 ;
    END
  END analog_io[23]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1387.325000 0.800000 1387.625000 ;
    END
  END analog_io[22]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1555.475000 0.800000 1555.775000 ;
    END
  END analog_io[21]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1723.625000 0.800000 1723.925000 ;
    END
  END analog_io[20]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1891.775000 0.800000 1892.075000 ;
    END
  END analog_io[19]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2059.925000 0.800000 2060.225000 ;
    END
  END analog_io[18]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2226.175000 0.800000 2226.475000 ;
    END
  END analog_io[17]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.630000 2289.750000 201.770000 2290.240000 ;
    END
  END analog_io[16]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.730000 2289.750000 470.870000 2290.240000 ;
    END
  END analog_io[15]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 739.830000 2289.750000 739.970000 2290.240000 ;
    END
  END analog_io[14]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1009.130000 2289.750000 1009.270000 2290.240000 ;
    END
  END analog_io[13]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1278.230000 2289.750000 1278.370000 2290.240000 ;
    END
  END analog_io[12]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1547.330000 2289.750000 1547.470000 2290.240000 ;
    END
  END analog_io[11]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1816.430000 2289.750000 1816.570000 2290.240000 ;
    END
  END analog_io[10]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2085.630000 2289.750000 2085.770000 2290.240000 ;
    END
  END analog_io[9]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2350.030000 2289.755000 2350.170000 2290.240000 ;
    END
  END analog_io[8]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 2099.635000 2369.460000 2099.935000 ;
    END
  END analog_io[7]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 1928.255000 2369.460000 1928.555000 ;
    END
  END analog_io[6]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 1756.780000 2369.460000 1757.080000 ;
    END
  END analog_io[5]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 1585.305000 2369.460000 1585.605000 ;
    END
  END analog_io[4]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 1413.925000 2369.460000 1414.225000 ;
    END
  END analog_io[3]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 1242.640000 2369.460000 1242.940000 ;
    END
  END analog_io[2]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 1071.070000 2369.460000 1071.370000 ;
    END
  END analog_io[1]
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2368.660000 899.690000 2369.460000 899.990000 ;
    END
  END analog_io[0]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2339.930000 0.000000 2340.070000 0.490000 ;
    END
  END user_clock2
  PIN user_irq[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9399 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.5915 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2356.730000 0.000000 2356.870000 0.485000 ;
    END
  END user_irq[2]
  PIN user_irq[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4236 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.01 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2349.430000 0.000000 2349.570000 0.490000 ;
    END
  END user_irq[1]
  PIN user_irq[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9154 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.469 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2344.630000 0.000000 2344.770000 0.490000 ;
    END
  END user_irq[0]
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 7.980000 8.260000 2361.480000 12.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.980000 2277.300000 2361.480000 2281.300000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2357.480000 8.260000 2361.480000 2281.300000 ;
    END
    PORT
      LAYER met4 ;
        RECT 7.980000 8.260000 11.980000 2281.300000 ;
    END

# P/G pin shape extracted from block 'tcam_32x28'
    PORT
      LAYER met4 ;
        RECT 668.435000 1811.260000 670.175000 2206.040000 ;
      LAYER met3 ;
        RECT 668.435000 2204.300000 1145.495000 2206.040000 ;
      LAYER met3 ;
        RECT 668.435000 1811.260000 1145.495000 1813.000000 ;
      LAYER met4 ;
        RECT 1143.755000 1811.260000 1145.495000 2206.040000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1230.575000 1811.355000 1232.315000 2206.135000 ;
      LAYER met3 ;
        RECT 1230.575000 2204.395000 1707.635000 2206.135000 ;
      LAYER met3 ;
        RECT 1230.575000 1811.355000 1707.635000 1813.095000 ;
      LAYER met4 ;
        RECT 1705.895000 1811.355000 1707.635000 2206.135000 ;
    END
    PORT
      LAYER met4 ;
        RECT 642.365000 1771.825000 644.365000 2241.665000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1731.905000 1771.825000 1733.905000 2241.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 642.365000 2239.665000 1733.905000 2241.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 642.365000 1771.825000 1733.905000 1773.825000 ;
    END
# end of P/G pin shape extracted from block 'tcam_32x28'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 513.045000 525.515000 514.785000 920.295000 ;
      LAYER met3 ;
        RECT 37.725000 525.515000 514.785000 527.255000 ;
      LAYER met3 ;
        RECT 37.725000 918.555000 514.785000 920.295000 ;
      LAYER met4 ;
        RECT 37.725000 525.515000 39.465000 920.295000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 513.045000 967.215000 514.785000 1361.995000 ;
      LAYER met3 ;
        RECT 37.725000 967.215000 514.785000 968.955000 ;
      LAYER met3 ;
        RECT 37.725000 1360.255000 514.785000 1361.995000 ;
      LAYER met4 ;
        RECT 37.725000 967.215000 39.465000 1361.995000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 513.045000 1408.915000 514.785000 1803.695000 ;
      LAYER met3 ;
        RECT 37.725000 1408.915000 514.785000 1410.655000 ;
      LAYER met3 ;
        RECT 37.725000 1801.955000 514.785000 1803.695000 ;
      LAYER met4 ;
        RECT 37.725000 1408.915000 39.465000 1803.695000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 513.045000 1850.615000 514.785000 2245.395000 ;
      LAYER met3 ;
        RECT 37.725000 1850.615000 514.785000 1852.355000 ;
      LAYER met3 ;
        RECT 37.725000 2243.655000 514.785000 2245.395000 ;
      LAYER met4 ;
        RECT 37.725000 1850.615000 39.465000 2245.395000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 2335.145000 525.515000 2336.885000 920.295000 ;
      LAYER met3 ;
        RECT 1859.825000 525.515000 2336.885000 527.255000 ;
      LAYER met3 ;
        RECT 1859.825000 918.555000 2336.885000 920.295000 ;
      LAYER met4 ;
        RECT 1859.825000 525.515000 1861.565000 920.295000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 2335.145000 967.215000 2336.885000 1361.995000 ;
      LAYER met3 ;
        RECT 1859.825000 967.215000 2336.885000 968.955000 ;
      LAYER met3 ;
        RECT 1859.825000 1360.255000 2336.885000 1361.995000 ;
      LAYER met4 ;
        RECT 1859.825000 967.215000 1861.565000 1361.995000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 2335.145000 1408.915000 2336.885000 1803.695000 ;
      LAYER met3 ;
        RECT 1859.825000 1408.915000 2336.885000 1410.655000 ;
      LAYER met3 ;
        RECT 1859.825000 1801.955000 2336.885000 1803.695000 ;
      LAYER met4 ;
        RECT 1859.825000 1408.915000 1861.565000 1803.695000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 2335.145000 1850.615000 2336.885000 2245.395000 ;
      LAYER met3 ;
        RECT 1859.825000 1850.615000 2336.885000 1852.355000 ;
      LAYER met3 ;
        RECT 1859.825000 2243.655000 2336.885000 2245.395000 ;
      LAYER met4 ;
        RECT 1859.825000 1850.615000 1861.565000 2245.395000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END vssd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 13.780000 14.060000 2355.680000 18.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780000 2271.500000 2355.680000 2275.500000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2351.680000 14.060000 2355.680000 2275.500000 ;
    END
    PORT
      LAYER met4 ;
        RECT 13.780000 14.060000 17.780000 2275.500000 ;
    END

# P/G pin shape extracted from block 'tcam_32x28'
    PORT
      LAYER met4 ;
        RECT 1140.355000 1814.660000 1142.095000 2202.640000 ;
      LAYER met4 ;
        RECT 671.835000 1814.660000 673.575000 2202.640000 ;
      LAYER met3 ;
        RECT 671.835000 1814.660000 1142.095000 1816.400000 ;
      LAYER met3 ;
        RECT 671.835000 2200.900000 1142.095000 2202.640000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1702.495000 1814.755000 1704.235000 2202.735000 ;
      LAYER met4 ;
        RECT 1233.975000 1814.755000 1235.715000 2202.735000 ;
      LAYER met3 ;
        RECT 1233.975000 1814.755000 1704.235000 1816.495000 ;
      LAYER met3 ;
        RECT 1233.975000 2200.995000 1704.235000 2202.735000 ;
    END
    PORT
      LAYER met4 ;
        RECT 646.165000 1775.625000 648.165000 2237.865000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1728.105000 1775.625000 1730.105000 2237.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 646.165000 2235.865000 1730.105000 2237.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 646.165000 1775.625000 1730.105000 1777.625000 ;
    END
# end of P/G pin shape extracted from block 'tcam_32x28'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 41.125000 915.155000 511.385000 916.895000 ;
      LAYER met3 ;
        RECT 41.125000 528.915000 511.385000 530.655000 ;
      LAYER met4 ;
        RECT 41.125000 528.915000 42.865000 916.895000 ;
      LAYER met4 ;
        RECT 509.645000 528.915000 511.385000 916.895000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 41.125000 1356.855000 511.385000 1358.595000 ;
      LAYER met3 ;
        RECT 41.125000 970.615000 511.385000 972.355000 ;
      LAYER met4 ;
        RECT 41.125000 970.615000 42.865000 1358.595000 ;
      LAYER met4 ;
        RECT 509.645000 970.615000 511.385000 1358.595000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 41.125000 1798.555000 511.385000 1800.295000 ;
      LAYER met3 ;
        RECT 41.125000 1412.315000 511.385000 1414.055000 ;
      LAYER met4 ;
        RECT 41.125000 1412.315000 42.865000 1800.295000 ;
      LAYER met4 ;
        RECT 509.645000 1412.315000 511.385000 1800.295000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 41.125000 2240.255000 511.385000 2241.995000 ;
      LAYER met3 ;
        RECT 41.125000 1854.015000 511.385000 1855.755000 ;
      LAYER met4 ;
        RECT 41.125000 1854.015000 42.865000 2241.995000 ;
      LAYER met4 ;
        RECT 509.645000 1854.015000 511.385000 2241.995000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 1863.225000 915.155000 2333.485000 916.895000 ;
      LAYER met3 ;
        RECT 1863.225000 528.915000 2333.485000 530.655000 ;
      LAYER met4 ;
        RECT 1863.225000 528.915000 1864.965000 916.895000 ;
      LAYER met4 ;
        RECT 2331.745000 528.915000 2333.485000 916.895000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 1863.225000 1356.855000 2333.485000 1358.595000 ;
      LAYER met3 ;
        RECT 1863.225000 970.615000 2333.485000 972.355000 ;
      LAYER met4 ;
        RECT 1863.225000 970.615000 1864.965000 1358.595000 ;
      LAYER met4 ;
        RECT 2331.745000 970.615000 2333.485000 1358.595000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 1863.225000 1798.555000 2333.485000 1800.295000 ;
      LAYER met3 ;
        RECT 1863.225000 1412.315000 2333.485000 1414.055000 ;
      LAYER met4 ;
        RECT 1863.225000 1412.315000 1864.965000 1800.295000 ;
      LAYER met4 ;
        RECT 2331.745000 1412.315000 2333.485000 1800.295000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 1863.225000 2240.255000 2333.485000 2241.995000 ;
      LAYER met3 ;
        RECT 1863.225000 1854.015000 2333.485000 1855.755000 ;
      LAYER met4 ;
        RECT 1863.225000 1854.015000 1864.965000 2241.995000 ;
      LAYER met4 ;
        RECT 2331.745000 1854.015000 2333.485000 2241.995000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END vccd1
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 2369.460000 2290.240000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 2369.460000 2290.240000 ;
    LAYER met2 ;
      RECT 2350.310000 2289.615000 2369.460000 2290.240000 ;
      RECT 2287.710000 2289.615000 2349.890000 2290.240000 ;
      RECT 5.010000 2289.615000 66.890000 2290.240000 ;
      RECT 0.000000 2289.615000 4.590000 2290.240000 ;
      RECT 2287.710000 2289.610000 2369.460000 2289.615000 ;
      RECT 2220.310000 2289.610000 2287.290000 2290.240000 ;
      RECT 2153.110000 2289.610000 2219.890000 2290.240000 ;
      RECT 2085.910000 2289.610000 2152.690000 2290.240000 ;
      RECT 2018.610000 2289.610000 2085.490000 2290.240000 ;
      RECT 1951.210000 2289.610000 2018.190000 2290.240000 ;
      RECT 1884.010000 2289.610000 1950.790000 2290.240000 ;
      RECT 1816.710000 2289.610000 1883.590000 2290.240000 ;
      RECT 1749.410000 2289.610000 1816.290000 2290.240000 ;
      RECT 1682.110000 2289.610000 1748.990000 2290.240000 ;
      RECT 1614.910000 2289.610000 1681.690000 2290.240000 ;
      RECT 1547.610000 2289.610000 1614.490000 2290.240000 ;
      RECT 1480.310000 2289.610000 1547.190000 2290.240000 ;
      RECT 1413.010000 2289.610000 1479.890000 2290.240000 ;
      RECT 1345.710000 2289.610000 1412.590000 2290.240000 ;
      RECT 1278.510000 2289.610000 1345.290000 2290.240000 ;
      RECT 1211.110000 2289.610000 1278.090000 2290.240000 ;
      RECT 1143.810000 2289.610000 1210.690000 2290.240000 ;
      RECT 1076.610000 2289.610000 1143.390000 2290.240000 ;
      RECT 1009.410000 2289.610000 1076.190000 2290.240000 ;
      RECT 942.010000 2289.610000 1008.990000 2290.240000 ;
      RECT 874.710000 2289.610000 941.590000 2290.240000 ;
      RECT 807.510000 2289.610000 874.290000 2290.240000 ;
      RECT 740.110000 2289.610000 807.090000 2290.240000 ;
      RECT 672.810000 2289.610000 739.690000 2290.240000 ;
      RECT 605.610000 2289.610000 672.390000 2290.240000 ;
      RECT 538.410000 2289.610000 605.190000 2290.240000 ;
      RECT 471.010000 2289.610000 537.990000 2290.240000 ;
      RECT 403.810000 2289.610000 470.590000 2290.240000 ;
      RECT 336.510000 2289.610000 403.390000 2290.240000 ;
      RECT 269.210000 2289.610000 336.090000 2290.240000 ;
      RECT 201.910000 2289.610000 268.790000 2290.240000 ;
      RECT 134.610000 2289.610000 201.490000 2290.240000 ;
      RECT 67.310000 2289.610000 134.190000 2290.240000 ;
      RECT 0.000000 2289.610000 66.890000 2289.615000 ;
      RECT 0.000000 0.630000 2369.460000 2289.610000 ;
      RECT 2349.710000 0.625000 2369.460000 0.630000 ;
      RECT 0.000000 0.625000 4.390000 0.630000 ;
      RECT 2357.010000 0.000000 2369.460000 0.625000 ;
      RECT 2349.710000 0.000000 2356.590000 0.625000 ;
      RECT 2344.910000 0.000000 2349.290000 0.630000 ;
      RECT 2340.210000 0.000000 2344.490000 0.630000 ;
      RECT 2335.410000 0.000000 2339.790000 0.630000 ;
      RECT 2330.610000 0.000000 2334.990000 0.630000 ;
      RECT 2325.810000 0.000000 2330.190000 0.630000 ;
      RECT 2321.010000 0.000000 2325.390000 0.630000 ;
      RECT 2316.210000 0.000000 2320.590000 0.630000 ;
      RECT 2311.410000 0.000000 2315.790000 0.630000 ;
      RECT 2306.710000 0.000000 2310.990000 0.630000 ;
      RECT 2302.010000 0.000000 2306.290000 0.630000 ;
      RECT 2297.210000 0.000000 2301.590000 0.630000 ;
      RECT 2292.410000 0.000000 2296.790000 0.630000 ;
      RECT 2287.610000 0.000000 2291.990000 0.630000 ;
      RECT 2282.810000 0.000000 2287.190000 0.630000 ;
      RECT 2278.110000 0.000000 2282.390000 0.630000 ;
      RECT 2273.310000 0.000000 2277.690000 0.630000 ;
      RECT 2268.510000 0.000000 2272.890000 0.630000 ;
      RECT 2263.710000 0.000000 2268.090000 0.630000 ;
      RECT 2258.910000 0.000000 2263.290000 0.630000 ;
      RECT 2254.210000 0.000000 2258.490000 0.630000 ;
      RECT 2249.510000 0.000000 2253.790000 0.630000 ;
      RECT 2244.710000 0.000000 2249.090000 0.630000 ;
      RECT 2239.910000 0.000000 2244.290000 0.630000 ;
      RECT 2235.110000 0.000000 2239.490000 0.630000 ;
      RECT 2230.310000 0.000000 2234.690000 0.630000 ;
      RECT 2225.510000 0.000000 2229.890000 0.630000 ;
      RECT 2220.810000 0.000000 2225.090000 0.630000 ;
      RECT 2216.010000 0.000000 2220.390000 0.630000 ;
      RECT 2211.210000 0.000000 2215.590000 0.630000 ;
      RECT 2206.510000 0.000000 2210.790000 0.630000 ;
      RECT 2201.710000 0.000000 2206.090000 0.630000 ;
      RECT 2196.910000 0.000000 2201.290000 0.630000 ;
      RECT 2192.210000 0.000000 2196.490000 0.630000 ;
      RECT 2187.410000 0.000000 2191.790000 0.630000 ;
      RECT 2182.610000 0.000000 2186.990000 0.630000 ;
      RECT 2177.810000 0.000000 2182.190000 0.630000 ;
      RECT 2173.010000 0.000000 2177.390000 0.630000 ;
      RECT 2168.210000 0.000000 2172.590000 0.630000 ;
      RECT 2163.510000 0.000000 2167.790000 0.630000 ;
      RECT 2158.810000 0.000000 2163.090000 0.630000 ;
      RECT 2154.010000 0.000000 2158.390000 0.630000 ;
      RECT 2149.210000 0.000000 2153.590000 0.630000 ;
      RECT 2144.410000 0.000000 2148.790000 0.630000 ;
      RECT 2139.510000 0.000000 2143.990000 0.630000 ;
      RECT 2134.810000 0.000000 2139.090000 0.630000 ;
      RECT 2130.010000 0.000000 2134.390000 0.630000 ;
      RECT 2125.210000 0.000000 2129.590000 0.630000 ;
      RECT 2120.410000 0.000000 2124.790000 0.630000 ;
      RECT 2115.610000 0.000000 2119.990000 0.630000 ;
      RECT 2110.810000 0.000000 2115.190000 0.630000 ;
      RECT 2106.210000 0.000000 2110.390000 0.630000 ;
      RECT 2101.410000 0.000000 2105.790000 0.630000 ;
      RECT 2096.610000 0.000000 2100.990000 0.630000 ;
      RECT 2091.810000 0.000000 2096.190000 0.630000 ;
      RECT 2087.010000 0.000000 2091.390000 0.630000 ;
      RECT 2082.210000 0.000000 2086.590000 0.630000 ;
      RECT 2077.410000 0.000000 2081.790000 0.630000 ;
      RECT 2072.710000 0.000000 2076.990000 0.630000 ;
      RECT 2067.910000 0.000000 2072.290000 0.630000 ;
      RECT 2063.110000 0.000000 2067.490000 0.630000 ;
      RECT 2058.410000 0.000000 2062.690000 0.630000 ;
      RECT 2053.610000 0.000000 2057.990000 0.630000 ;
      RECT 2048.810000 0.000000 2053.190000 0.630000 ;
      RECT 2044.110000 0.000000 2048.390000 0.630000 ;
      RECT 2039.310000 0.000000 2043.690000 0.630000 ;
      RECT 2034.510000 0.000000 2038.890000 0.630000 ;
      RECT 2029.710000 0.000000 2034.090000 0.630000 ;
      RECT 2024.910000 0.000000 2029.290000 0.630000 ;
      RECT 2020.110000 0.000000 2024.490000 0.630000 ;
      RECT 2015.410000 0.000000 2019.690000 0.630000 ;
      RECT 2010.710000 0.000000 2014.990000 0.630000 ;
      RECT 2005.910000 0.000000 2010.290000 0.630000 ;
      RECT 2001.110000 0.000000 2005.490000 0.630000 ;
      RECT 1996.310000 0.000000 2000.690000 0.630000 ;
      RECT 1991.510000 0.000000 1995.890000 0.630000 ;
      RECT 1986.810000 0.000000 1991.090000 0.630000 ;
      RECT 1982.010000 0.000000 1986.390000 0.630000 ;
      RECT 1977.210000 0.000000 1981.590000 0.630000 ;
      RECT 1972.410000 0.000000 1976.790000 0.630000 ;
      RECT 1967.610000 0.000000 1971.990000 0.630000 ;
      RECT 1962.910000 0.000000 1967.190000 0.630000 ;
      RECT 1958.210000 0.000000 1962.490000 0.630000 ;
      RECT 1953.410000 0.000000 1957.790000 0.630000 ;
      RECT 1948.610000 0.000000 1952.990000 0.630000 ;
      RECT 1943.810000 0.000000 1948.190000 0.630000 ;
      RECT 1939.010000 0.000000 1943.390000 0.630000 ;
      RECT 1934.210000 0.000000 1938.590000 0.630000 ;
      RECT 1929.510000 0.000000 1933.790000 0.630000 ;
      RECT 1924.710000 0.000000 1929.090000 0.630000 ;
      RECT 1919.910000 0.000000 1924.290000 0.630000 ;
      RECT 1915.210000 0.000000 1919.490000 0.630000 ;
      RECT 1910.410000 0.000000 1914.790000 0.630000 ;
      RECT 1905.610000 0.000000 1909.990000 0.630000 ;
      RECT 1900.810000 0.000000 1905.190000 0.630000 ;
      RECT 1896.010000 0.000000 1900.390000 0.630000 ;
      RECT 1891.210000 0.000000 1895.590000 0.630000 ;
      RECT 1886.410000 0.000000 1890.790000 0.630000 ;
      RECT 1881.610000 0.000000 1885.990000 0.630000 ;
      RECT 1876.810000 0.000000 1881.190000 0.630000 ;
      RECT 1872.010000 0.000000 1876.390000 0.630000 ;
      RECT 1867.410000 0.000000 1871.590000 0.630000 ;
      RECT 1862.610000 0.000000 1866.990000 0.630000 ;
      RECT 1857.810000 0.000000 1862.190000 0.630000 ;
      RECT 1853.010000 0.000000 1857.390000 0.630000 ;
      RECT 1848.210000 0.000000 1852.590000 0.630000 ;
      RECT 1843.410000 0.000000 1847.790000 0.630000 ;
      RECT 1838.710000 0.000000 1842.990000 0.630000 ;
      RECT 1833.910000 0.000000 1838.290000 0.630000 ;
      RECT 1829.110000 0.000000 1833.490000 0.630000 ;
      RECT 1824.310000 0.000000 1828.690000 0.630000 ;
      RECT 1819.610000 0.000000 1823.890000 0.630000 ;
      RECT 1814.810000 0.000000 1819.190000 0.630000 ;
      RECT 1810.110000 0.000000 1814.390000 0.630000 ;
      RECT 1805.310000 0.000000 1809.690000 0.630000 ;
      RECT 1800.510000 0.000000 1804.890000 0.630000 ;
      RECT 1795.710000 0.000000 1800.090000 0.630000 ;
      RECT 1790.910000 0.000000 1795.290000 0.630000 ;
      RECT 1786.110000 0.000000 1790.490000 0.630000 ;
      RECT 1781.410000 0.000000 1785.690000 0.630000 ;
      RECT 1776.610000 0.000000 1780.990000 0.630000 ;
      RECT 1771.910000 0.000000 1776.190000 0.630000 ;
      RECT 1767.110000 0.000000 1771.490000 0.630000 ;
      RECT 1762.310000 0.000000 1766.690000 0.630000 ;
      RECT 1757.510000 0.000000 1761.890000 0.630000 ;
      RECT 1752.810000 0.000000 1757.090000 0.630000 ;
      RECT 1748.010000 0.000000 1752.390000 0.630000 ;
      RECT 1743.210000 0.000000 1747.590000 0.630000 ;
      RECT 1738.410000 0.000000 1742.790000 0.630000 ;
      RECT 1733.610000 0.000000 1737.990000 0.630000 ;
      RECT 1728.810000 0.000000 1733.190000 0.630000 ;
      RECT 1724.210000 0.000000 1728.390000 0.630000 ;
      RECT 1719.410000 0.000000 1723.790000 0.630000 ;
      RECT 1714.610000 0.000000 1718.990000 0.630000 ;
      RECT 1709.810000 0.000000 1714.190000 0.630000 ;
      RECT 1705.010000 0.000000 1709.390000 0.630000 ;
      RECT 1700.210000 0.000000 1704.590000 0.630000 ;
      RECT 1695.510000 0.000000 1699.790000 0.630000 ;
      RECT 1690.710000 0.000000 1695.090000 0.630000 ;
      RECT 1685.910000 0.000000 1690.290000 0.630000 ;
      RECT 1681.110000 0.000000 1685.490000 0.630000 ;
      RECT 1676.410000 0.000000 1680.690000 0.630000 ;
      RECT 1671.610000 0.000000 1675.990000 0.630000 ;
      RECT 1666.910000 0.000000 1671.190000 0.630000 ;
      RECT 1662.010000 0.000000 1666.490000 0.630000 ;
      RECT 1657.210000 0.000000 1661.590000 0.630000 ;
      RECT 1652.410000 0.000000 1656.790000 0.630000 ;
      RECT 1647.610000 0.000000 1651.990000 0.630000 ;
      RECT 1642.810000 0.000000 1647.190000 0.630000 ;
      RECT 1638.010000 0.000000 1642.390000 0.630000 ;
      RECT 1633.310000 0.000000 1637.590000 0.630000 ;
      RECT 1628.610000 0.000000 1632.890000 0.630000 ;
      RECT 1623.810000 0.000000 1628.190000 0.630000 ;
      RECT 1619.010000 0.000000 1623.390000 0.630000 ;
      RECT 1614.210000 0.000000 1618.590000 0.630000 ;
      RECT 1609.410000 0.000000 1613.790000 0.630000 ;
      RECT 1604.710000 0.000000 1608.990000 0.630000 ;
      RECT 1599.910000 0.000000 1604.290000 0.630000 ;
      RECT 1595.110000 0.000000 1599.490000 0.630000 ;
      RECT 1590.310000 0.000000 1594.690000 0.630000 ;
      RECT 1585.510000 0.000000 1589.890000 0.630000 ;
      RECT 1580.810000 0.000000 1585.090000 0.630000 ;
      RECT 1576.110000 0.000000 1580.390000 0.630000 ;
      RECT 1571.310000 0.000000 1575.690000 0.630000 ;
      RECT 1566.510000 0.000000 1570.890000 0.630000 ;
      RECT 1561.710000 0.000000 1566.090000 0.630000 ;
      RECT 1556.910000 0.000000 1561.290000 0.630000 ;
      RECT 1552.110000 0.000000 1556.490000 0.630000 ;
      RECT 1547.410000 0.000000 1551.690000 0.630000 ;
      RECT 1542.610000 0.000000 1546.990000 0.630000 ;
      RECT 1537.810000 0.000000 1542.190000 0.630000 ;
      RECT 1533.110000 0.000000 1537.390000 0.630000 ;
      RECT 1528.310000 0.000000 1532.690000 0.630000 ;
      RECT 1523.510000 0.000000 1527.890000 0.630000 ;
      RECT 1518.810000 0.000000 1523.090000 0.630000 ;
      RECT 1514.010000 0.000000 1518.390000 0.630000 ;
      RECT 1509.210000 0.000000 1513.590000 0.630000 ;
      RECT 1504.410000 0.000000 1508.790000 0.630000 ;
      RECT 1499.610000 0.000000 1503.990000 0.630000 ;
      RECT 1494.810000 0.000000 1499.190000 0.630000 ;
      RECT 1490.110000 0.000000 1494.390000 0.630000 ;
      RECT 1485.410000 0.000000 1489.690000 0.630000 ;
      RECT 1480.610000 0.000000 1484.990000 0.630000 ;
      RECT 1475.810000 0.000000 1480.190000 0.630000 ;
      RECT 1471.010000 0.000000 1475.390000 0.630000 ;
      RECT 1466.210000 0.000000 1470.590000 0.630000 ;
      RECT 1461.510000 0.000000 1465.790000 0.630000 ;
      RECT 1456.710000 0.000000 1461.090000 0.630000 ;
      RECT 1451.910000 0.000000 1456.290000 0.630000 ;
      RECT 1447.110000 0.000000 1451.490000 0.630000 ;
      RECT 1442.310000 0.000000 1446.690000 0.630000 ;
      RECT 1437.610000 0.000000 1441.890000 0.630000 ;
      RECT 1432.910000 0.000000 1437.190000 0.630000 ;
      RECT 1428.110000 0.000000 1432.490000 0.630000 ;
      RECT 1423.210000 0.000000 1427.690000 0.630000 ;
      RECT 1418.410000 0.000000 1422.790000 0.630000 ;
      RECT 1413.610000 0.000000 1417.990000 0.630000 ;
      RECT 1408.810000 0.000000 1413.190000 0.630000 ;
      RECT 1404.010000 0.000000 1408.390000 0.630000 ;
      RECT 1399.310000 0.000000 1403.590000 0.630000 ;
      RECT 1394.510000 0.000000 1398.890000 0.630000 ;
      RECT 1389.810000 0.000000 1394.090000 0.630000 ;
      RECT 1385.010000 0.000000 1389.390000 0.630000 ;
      RECT 1380.210000 0.000000 1384.590000 0.630000 ;
      RECT 1375.410000 0.000000 1379.790000 0.630000 ;
      RECT 1370.710000 0.000000 1374.990000 0.630000 ;
      RECT 1365.910000 0.000000 1370.290000 0.630000 ;
      RECT 1361.110000 0.000000 1365.490000 0.630000 ;
      RECT 1356.310000 0.000000 1360.690000 0.630000 ;
      RECT 1351.510000 0.000000 1355.890000 0.630000 ;
      RECT 1346.710000 0.000000 1351.090000 0.630000 ;
      RECT 1342.110000 0.000000 1346.290000 0.630000 ;
      RECT 1337.310000 0.000000 1341.690000 0.630000 ;
      RECT 1332.510000 0.000000 1336.890000 0.630000 ;
      RECT 1327.710000 0.000000 1332.090000 0.630000 ;
      RECT 1322.910000 0.000000 1327.290000 0.630000 ;
      RECT 1318.110000 0.000000 1322.490000 0.630000 ;
      RECT 1313.410000 0.000000 1317.690000 0.630000 ;
      RECT 1308.610000 0.000000 1312.990000 0.630000 ;
      RECT 1303.810000 0.000000 1308.190000 0.630000 ;
      RECT 1299.010000 0.000000 1303.390000 0.630000 ;
      RECT 1294.310000 0.000000 1298.590000 0.630000 ;
      RECT 1289.510000 0.000000 1293.890000 0.630000 ;
      RECT 1284.810000 0.000000 1289.090000 0.630000 ;
      RECT 1280.010000 0.000000 1284.390000 0.630000 ;
      RECT 1275.210000 0.000000 1279.590000 0.630000 ;
      RECT 1270.410000 0.000000 1274.790000 0.630000 ;
      RECT 1265.610000 0.000000 1269.990000 0.630000 ;
      RECT 1260.810000 0.000000 1265.190000 0.630000 ;
      RECT 1256.110000 0.000000 1260.390000 0.630000 ;
      RECT 1251.310000 0.000000 1255.690000 0.630000 ;
      RECT 1246.610000 0.000000 1250.890000 0.630000 ;
      RECT 1241.810000 0.000000 1246.190000 0.630000 ;
      RECT 1237.010000 0.000000 1241.390000 0.630000 ;
      RECT 1232.210000 0.000000 1236.590000 0.630000 ;
      RECT 1227.510000 0.000000 1231.790000 0.630000 ;
      RECT 1222.710000 0.000000 1227.090000 0.630000 ;
      RECT 1217.910000 0.000000 1222.290000 0.630000 ;
      RECT 1213.110000 0.000000 1217.490000 0.630000 ;
      RECT 1208.310000 0.000000 1212.690000 0.630000 ;
      RECT 1203.510000 0.000000 1207.890000 0.630000 ;
      RECT 1198.910000 0.000000 1203.090000 0.630000 ;
      RECT 1194.110000 0.000000 1198.490000 0.630000 ;
      RECT 1189.310000 0.000000 1193.690000 0.630000 ;
      RECT 1184.410000 0.000000 1188.890000 0.630000 ;
      RECT 1179.610000 0.000000 1183.990000 0.630000 ;
      RECT 1174.810000 0.000000 1179.190000 0.630000 ;
      RECT 1170.010000 0.000000 1174.390000 0.630000 ;
      RECT 1165.310000 0.000000 1169.590000 0.630000 ;
      RECT 1160.510000 0.000000 1164.890000 0.630000 ;
      RECT 1155.710000 0.000000 1160.090000 0.630000 ;
      RECT 1151.010000 0.000000 1155.290000 0.630000 ;
      RECT 1146.210000 0.000000 1150.590000 0.630000 ;
      RECT 1141.410000 0.000000 1145.790000 0.630000 ;
      RECT 1136.710000 0.000000 1140.990000 0.630000 ;
      RECT 1131.910000 0.000000 1136.290000 0.630000 ;
      RECT 1127.110000 0.000000 1131.490000 0.630000 ;
      RECT 1122.310000 0.000000 1126.690000 0.630000 ;
      RECT 1117.510000 0.000000 1121.890000 0.630000 ;
      RECT 1112.710000 0.000000 1117.090000 0.630000 ;
      RECT 1108.010000 0.000000 1112.290000 0.630000 ;
      RECT 1103.310000 0.000000 1107.590000 0.630000 ;
      RECT 1098.510000 0.000000 1102.890000 0.630000 ;
      RECT 1093.710000 0.000000 1098.090000 0.630000 ;
      RECT 1088.910000 0.000000 1093.290000 0.630000 ;
      RECT 1084.110000 0.000000 1088.490000 0.630000 ;
      RECT 1079.410000 0.000000 1083.690000 0.630000 ;
      RECT 1074.610000 0.000000 1078.990000 0.630000 ;
      RECT 1069.810000 0.000000 1074.190000 0.630000 ;
      RECT 1065.010000 0.000000 1069.390000 0.630000 ;
      RECT 1060.210000 0.000000 1064.590000 0.630000 ;
      RECT 1055.510000 0.000000 1059.790000 0.630000 ;
      RECT 1050.810000 0.000000 1055.090000 0.630000 ;
      RECT 1046.010000 0.000000 1050.390000 0.630000 ;
      RECT 1041.210000 0.000000 1045.590000 0.630000 ;
      RECT 1036.410000 0.000000 1040.790000 0.630000 ;
      RECT 1031.610000 0.000000 1035.990000 0.630000 ;
      RECT 1026.810000 0.000000 1031.190000 0.630000 ;
      RECT 1022.110000 0.000000 1026.390000 0.630000 ;
      RECT 1017.310000 0.000000 1021.690000 0.630000 ;
      RECT 1012.510000 0.000000 1016.890000 0.630000 ;
      RECT 1007.810000 0.000000 1012.090000 0.630000 ;
      RECT 1003.010000 0.000000 1007.390000 0.630000 ;
      RECT 998.210000 0.000000 1002.590000 0.630000 ;
      RECT 993.510000 0.000000 997.790000 0.630000 ;
      RECT 988.710000 0.000000 993.090000 0.630000 ;
      RECT 983.910000 0.000000 988.290000 0.630000 ;
      RECT 979.110000 0.000000 983.490000 0.630000 ;
      RECT 974.310000 0.000000 978.690000 0.630000 ;
      RECT 969.510000 0.000000 973.890000 0.630000 ;
      RECT 964.810000 0.000000 969.090000 0.630000 ;
      RECT 960.110000 0.000000 964.390000 0.630000 ;
      RECT 955.310000 0.000000 959.690000 0.630000 ;
      RECT 950.510000 0.000000 954.890000 0.630000 ;
      RECT 945.610000 0.000000 950.090000 0.630000 ;
      RECT 940.810000 0.000000 945.190000 0.630000 ;
      RECT 936.010000 0.000000 940.390000 0.630000 ;
      RECT 931.310000 0.000000 935.590000 0.630000 ;
      RECT 926.510000 0.000000 930.890000 0.630000 ;
      RECT 921.710000 0.000000 926.090000 0.630000 ;
      RECT 916.910000 0.000000 921.290000 0.630000 ;
      RECT 912.110000 0.000000 916.490000 0.630000 ;
      RECT 907.410000 0.000000 911.690000 0.630000 ;
      RECT 902.710000 0.000000 906.990000 0.630000 ;
      RECT 897.910000 0.000000 902.290000 0.630000 ;
      RECT 893.110000 0.000000 897.490000 0.630000 ;
      RECT 888.310000 0.000000 892.690000 0.630000 ;
      RECT 883.510000 0.000000 887.890000 0.630000 ;
      RECT 878.710000 0.000000 883.090000 0.630000 ;
      RECT 874.010000 0.000000 878.290000 0.630000 ;
      RECT 869.210000 0.000000 873.590000 0.630000 ;
      RECT 864.410000 0.000000 868.790000 0.630000 ;
      RECT 859.710000 0.000000 863.990000 0.630000 ;
      RECT 854.910000 0.000000 859.290000 0.630000 ;
      RECT 850.110000 0.000000 854.490000 0.630000 ;
      RECT 845.410000 0.000000 849.690000 0.630000 ;
      RECT 840.610000 0.000000 844.990000 0.630000 ;
      RECT 835.810000 0.000000 840.190000 0.630000 ;
      RECT 831.010000 0.000000 835.390000 0.630000 ;
      RECT 826.210000 0.000000 830.590000 0.630000 ;
      RECT 821.410000 0.000000 825.790000 0.630000 ;
      RECT 816.710000 0.000000 820.990000 0.630000 ;
      RECT 812.010000 0.000000 816.290000 0.630000 ;
      RECT 807.210000 0.000000 811.590000 0.630000 ;
      RECT 802.410000 0.000000 806.790000 0.630000 ;
      RECT 797.610000 0.000000 801.990000 0.630000 ;
      RECT 792.810000 0.000000 797.190000 0.630000 ;
      RECT 788.110000 0.000000 792.390000 0.630000 ;
      RECT 783.310000 0.000000 787.690000 0.630000 ;
      RECT 778.510000 0.000000 782.890000 0.630000 ;
      RECT 773.710000 0.000000 778.090000 0.630000 ;
      RECT 768.910000 0.000000 773.290000 0.630000 ;
      RECT 764.210000 0.000000 768.490000 0.630000 ;
      RECT 759.510000 0.000000 763.790000 0.630000 ;
      RECT 754.710000 0.000000 759.090000 0.630000 ;
      RECT 749.910000 0.000000 754.290000 0.630000 ;
      RECT 745.110000 0.000000 749.490000 0.630000 ;
      RECT 740.310000 0.000000 744.690000 0.630000 ;
      RECT 735.510000 0.000000 739.890000 0.630000 ;
      RECT 730.810000 0.000000 735.090000 0.630000 ;
      RECT 726.010000 0.000000 730.390000 0.630000 ;
      RECT 721.210000 0.000000 725.590000 0.630000 ;
      RECT 716.510000 0.000000 720.790000 0.630000 ;
      RECT 711.710000 0.000000 716.090000 0.630000 ;
      RECT 706.810000 0.000000 711.290000 0.630000 ;
      RECT 702.010000 0.000000 706.390000 0.630000 ;
      RECT 697.310000 0.000000 701.590000 0.630000 ;
      RECT 692.510000 0.000000 696.890000 0.630000 ;
      RECT 687.710000 0.000000 692.090000 0.630000 ;
      RECT 682.910000 0.000000 687.290000 0.630000 ;
      RECT 678.110000 0.000000 682.490000 0.630000 ;
      RECT 673.310000 0.000000 677.690000 0.630000 ;
      RECT 668.710000 0.000000 672.890000 0.630000 ;
      RECT 663.910000 0.000000 668.290000 0.630000 ;
      RECT 659.110000 0.000000 663.490000 0.630000 ;
      RECT 654.310000 0.000000 658.690000 0.630000 ;
      RECT 649.510000 0.000000 653.890000 0.630000 ;
      RECT 644.710000 0.000000 649.090000 0.630000 ;
      RECT 640.010000 0.000000 644.290000 0.630000 ;
      RECT 635.210000 0.000000 639.590000 0.630000 ;
      RECT 630.410000 0.000000 634.790000 0.630000 ;
      RECT 625.610000 0.000000 629.990000 0.630000 ;
      RECT 620.910000 0.000000 625.190000 0.630000 ;
      RECT 616.110000 0.000000 620.490000 0.630000 ;
      RECT 611.410000 0.000000 615.690000 0.630000 ;
      RECT 606.610000 0.000000 610.990000 0.630000 ;
      RECT 601.810000 0.000000 606.190000 0.630000 ;
      RECT 597.010000 0.000000 601.390000 0.630000 ;
      RECT 592.210000 0.000000 596.590000 0.630000 ;
      RECT 587.410000 0.000000 591.790000 0.630000 ;
      RECT 582.710000 0.000000 586.990000 0.630000 ;
      RECT 577.910000 0.000000 582.290000 0.630000 ;
      RECT 573.210000 0.000000 577.490000 0.630000 ;
      RECT 568.410000 0.000000 572.790000 0.630000 ;
      RECT 563.610000 0.000000 567.990000 0.630000 ;
      RECT 558.810000 0.000000 563.190000 0.630000 ;
      RECT 554.110000 0.000000 558.390000 0.630000 ;
      RECT 549.310000 0.000000 553.690000 0.630000 ;
      RECT 544.510000 0.000000 548.890000 0.630000 ;
      RECT 539.710000 0.000000 544.090000 0.630000 ;
      RECT 534.910000 0.000000 539.290000 0.630000 ;
      RECT 530.110000 0.000000 534.490000 0.630000 ;
      RECT 525.510000 0.000000 529.690000 0.630000 ;
      RECT 520.710000 0.000000 525.090000 0.630000 ;
      RECT 515.910000 0.000000 520.290000 0.630000 ;
      RECT 511.110000 0.000000 515.490000 0.630000 ;
      RECT 506.310000 0.000000 510.690000 0.630000 ;
      RECT 501.510000 0.000000 505.890000 0.630000 ;
      RECT 496.810000 0.000000 501.090000 0.630000 ;
      RECT 492.010000 0.000000 496.390000 0.630000 ;
      RECT 487.210000 0.000000 491.590000 0.630000 ;
      RECT 482.410000 0.000000 486.790000 0.630000 ;
      RECT 477.710000 0.000000 481.990000 0.630000 ;
      RECT 472.910000 0.000000 477.290000 0.630000 ;
      RECT 468.010000 0.000000 472.490000 0.630000 ;
      RECT 463.310000 0.000000 467.590000 0.630000 ;
      RECT 458.510000 0.000000 462.890000 0.630000 ;
      RECT 453.710000 0.000000 458.090000 0.630000 ;
      RECT 448.910000 0.000000 453.290000 0.630000 ;
      RECT 444.110000 0.000000 448.490000 0.630000 ;
      RECT 439.310000 0.000000 443.690000 0.630000 ;
      RECT 434.610000 0.000000 438.890000 0.630000 ;
      RECT 429.910000 0.000000 434.190000 0.630000 ;
      RECT 425.110000 0.000000 429.490000 0.630000 ;
      RECT 420.310000 0.000000 424.690000 0.630000 ;
      RECT 415.510000 0.000000 419.890000 0.630000 ;
      RECT 410.710000 0.000000 415.090000 0.630000 ;
      RECT 406.010000 0.000000 410.290000 0.630000 ;
      RECT 401.210000 0.000000 405.590000 0.630000 ;
      RECT 396.410000 0.000000 400.790000 0.630000 ;
      RECT 391.610000 0.000000 395.990000 0.630000 ;
      RECT 386.810000 0.000000 391.190000 0.630000 ;
      RECT 382.110000 0.000000 386.390000 0.630000 ;
      RECT 377.410000 0.000000 381.690000 0.630000 ;
      RECT 372.610000 0.000000 376.990000 0.630000 ;
      RECT 367.810000 0.000000 372.190000 0.630000 ;
      RECT 363.010000 0.000000 367.390000 0.630000 ;
      RECT 358.210000 0.000000 362.590000 0.630000 ;
      RECT 353.410000 0.000000 357.790000 0.630000 ;
      RECT 348.710000 0.000000 352.990000 0.630000 ;
      RECT 343.910000 0.000000 348.290000 0.630000 ;
      RECT 339.110000 0.000000 343.490000 0.630000 ;
      RECT 334.410000 0.000000 338.690000 0.630000 ;
      RECT 329.610000 0.000000 333.990000 0.630000 ;
      RECT 324.810000 0.000000 329.190000 0.630000 ;
      RECT 320.110000 0.000000 324.390000 0.630000 ;
      RECT 315.310000 0.000000 319.690000 0.630000 ;
      RECT 310.510000 0.000000 314.890000 0.630000 ;
      RECT 305.710000 0.000000 310.090000 0.630000 ;
      RECT 300.910000 0.000000 305.290000 0.630000 ;
      RECT 296.110000 0.000000 300.490000 0.630000 ;
      RECT 291.410000 0.000000 295.690000 0.630000 ;
      RECT 286.710000 0.000000 290.990000 0.630000 ;
      RECT 281.910000 0.000000 286.290000 0.630000 ;
      RECT 277.110000 0.000000 281.490000 0.630000 ;
      RECT 272.310000 0.000000 276.690000 0.630000 ;
      RECT 267.510000 0.000000 271.890000 0.630000 ;
      RECT 262.810000 0.000000 267.090000 0.630000 ;
      RECT 258.010000 0.000000 262.390000 0.630000 ;
      RECT 253.210000 0.000000 257.590000 0.630000 ;
      RECT 248.410000 0.000000 252.790000 0.630000 ;
      RECT 243.610000 0.000000 247.990000 0.630000 ;
      RECT 238.910000 0.000000 243.190000 0.630000 ;
      RECT 234.210000 0.000000 238.490000 0.630000 ;
      RECT 229.310000 0.000000 233.790000 0.630000 ;
      RECT 224.510000 0.000000 228.890000 0.630000 ;
      RECT 219.710000 0.000000 224.090000 0.630000 ;
      RECT 214.910000 0.000000 219.290000 0.630000 ;
      RECT 210.110000 0.000000 214.490000 0.630000 ;
      RECT 205.310000 0.000000 209.690000 0.630000 ;
      RECT 200.610000 0.000000 204.890000 0.630000 ;
      RECT 195.810000 0.000000 200.190000 0.630000 ;
      RECT 191.110000 0.000000 195.390000 0.630000 ;
      RECT 186.310000 0.000000 190.690000 0.630000 ;
      RECT 181.510000 0.000000 185.890000 0.630000 ;
      RECT 176.710000 0.000000 181.090000 0.630000 ;
      RECT 172.010000 0.000000 176.290000 0.630000 ;
      RECT 167.210000 0.000000 171.590000 0.630000 ;
      RECT 162.410000 0.000000 166.790000 0.630000 ;
      RECT 157.610000 0.000000 161.990000 0.630000 ;
      RECT 152.810000 0.000000 157.190000 0.630000 ;
      RECT 148.010000 0.000000 152.390000 0.630000 ;
      RECT 143.410000 0.000000 147.590000 0.630000 ;
      RECT 138.610000 0.000000 142.990000 0.630000 ;
      RECT 133.810000 0.000000 138.190000 0.630000 ;
      RECT 129.010000 0.000000 133.390000 0.630000 ;
      RECT 124.210000 0.000000 128.590000 0.630000 ;
      RECT 119.410000 0.000000 123.790000 0.630000 ;
      RECT 114.710000 0.000000 118.990000 0.630000 ;
      RECT 109.910000 0.000000 114.290000 0.630000 ;
      RECT 105.110000 0.000000 109.490000 0.630000 ;
      RECT 100.310000 0.000000 104.690000 0.630000 ;
      RECT 95.610000 0.000000 99.890000 0.630000 ;
      RECT 90.810000 0.000000 95.190000 0.630000 ;
      RECT 86.110000 0.000000 90.390000 0.630000 ;
      RECT 81.310000 0.000000 85.690000 0.630000 ;
      RECT 76.510000 0.000000 80.890000 0.630000 ;
      RECT 71.710000 0.000000 76.090000 0.630000 ;
      RECT 66.910000 0.000000 71.290000 0.630000 ;
      RECT 62.110000 0.000000 66.490000 0.630000 ;
      RECT 57.410000 0.000000 61.690000 0.630000 ;
      RECT 52.610000 0.000000 56.990000 0.630000 ;
      RECT 47.910000 0.000000 52.190000 0.630000 ;
      RECT 43.110000 0.000000 47.490000 0.630000 ;
      RECT 38.310000 0.000000 42.690000 0.630000 ;
      RECT 33.510000 0.000000 37.890000 0.630000 ;
      RECT 28.810000 0.000000 33.090000 0.630000 ;
      RECT 24.010000 0.000000 28.390000 0.630000 ;
      RECT 19.210000 0.000000 23.590000 0.630000 ;
      RECT 14.410000 0.000000 18.790000 0.630000 ;
      RECT 9.610000 0.000000 13.990000 0.630000 ;
      RECT 4.810000 0.000000 9.190000 0.630000 ;
      RECT 2.210000 0.000000 4.390000 0.625000 ;
      RECT 0.000000 0.000000 1.790000 0.625000 ;
    LAYER met3 ;
      RECT 0.000000 2281.700000 2369.460000 2290.240000 ;
      RECT 2361.880000 2276.900000 2369.460000 2281.700000 ;
      RECT 0.000000 2276.900000 7.580000 2281.700000 ;
      RECT 0.000000 2275.900000 2369.460000 2276.900000 ;
      RECT 2356.080000 2271.100000 2369.460000 2275.900000 ;
      RECT 0.000000 2271.100000 13.380000 2275.900000 ;
      RECT 0.000000 2226.775000 2369.460000 2271.100000 ;
      RECT 1.100000 2225.875000 2369.460000 2226.775000 ;
      RECT 0.000000 2225.825000 2369.460000 2225.875000 ;
      RECT 0.000000 2224.925000 2368.360000 2225.825000 ;
      RECT 0.000000 2186.780000 2369.460000 2224.925000 ;
      RECT 1.100000 2186.020000 2369.460000 2186.780000 ;
      RECT 1.100000 2185.880000 2368.360000 2186.020000 ;
      RECT 0.000000 2185.120000 2368.360000 2185.880000 ;
      RECT 0.000000 2144.790000 2369.460000 2185.120000 ;
      RECT 1.100000 2143.890000 2369.460000 2144.790000 ;
      RECT 0.000000 2143.175000 2369.460000 2143.890000 ;
      RECT 0.000000 2142.275000 2368.360000 2143.175000 ;
      RECT 0.000000 2102.705000 2369.460000 2142.275000 ;
      RECT 1.100000 2101.805000 2369.460000 2102.705000 ;
      RECT 0.000000 2100.235000 2369.460000 2101.805000 ;
      RECT 0.000000 2099.335000 2368.360000 2100.235000 ;
      RECT 0.000000 2060.525000 2369.460000 2099.335000 ;
      RECT 1.100000 2059.625000 2369.460000 2060.525000 ;
      RECT 0.000000 2057.485000 2369.460000 2059.625000 ;
      RECT 0.000000 2056.585000 2368.360000 2057.485000 ;
      RECT 0.000000 2018.630000 2369.460000 2056.585000 ;
      RECT 1.100000 2017.730000 2369.460000 2018.630000 ;
      RECT 0.000000 2014.545000 2369.460000 2017.730000 ;
      RECT 0.000000 2013.645000 2368.360000 2014.545000 ;
      RECT 0.000000 1976.640000 2369.460000 2013.645000 ;
      RECT 1.100000 1975.740000 2369.460000 1976.640000 ;
      RECT 0.000000 1971.605000 2369.460000 1975.740000 ;
      RECT 0.000000 1970.705000 2368.360000 1971.605000 ;
      RECT 0.000000 1934.460000 2369.460000 1970.705000 ;
      RECT 1.100000 1933.560000 2369.460000 1934.460000 ;
      RECT 0.000000 1928.855000 2369.460000 1933.560000 ;
      RECT 0.000000 1927.955000 2368.360000 1928.855000 ;
      RECT 0.000000 1892.375000 2369.460000 1927.955000 ;
      RECT 1.100000 1891.475000 2369.460000 1892.375000 ;
      RECT 0.000000 1885.915000 2369.460000 1891.475000 ;
      RECT 0.000000 1885.015000 2368.360000 1885.915000 ;
      RECT 0.000000 1850.480000 2369.460000 1885.015000 ;
      RECT 1.100000 1849.580000 2369.460000 1850.480000 ;
      RECT 0.000000 1843.165000 2369.460000 1849.580000 ;
      RECT 0.000000 1842.265000 2368.360000 1843.165000 ;
      RECT 0.000000 1808.395000 2369.460000 1842.265000 ;
      RECT 1.100000 1807.495000 2369.460000 1808.395000 ;
      RECT 0.000000 1800.225000 2369.460000 1807.495000 ;
      RECT 0.000000 1799.325000 2368.360000 1800.225000 ;
      RECT 0.000000 1766.310000 2369.460000 1799.325000 ;
      RECT 1.100000 1765.410000 2369.460000 1766.310000 ;
      RECT 0.000000 1757.380000 2369.460000 1765.410000 ;
      RECT 0.000000 1756.480000 2368.360000 1757.380000 ;
      RECT 0.000000 1724.225000 2369.460000 1756.480000 ;
      RECT 1.100000 1723.325000 2369.460000 1724.225000 ;
      RECT 0.000000 1714.535000 2369.460000 1723.325000 ;
      RECT 0.000000 1713.635000 2368.360000 1714.535000 ;
      RECT 0.000000 1682.140000 2369.460000 1713.635000 ;
      RECT 1.100000 1681.240000 2369.460000 1682.140000 ;
      RECT 0.000000 1671.690000 2369.460000 1681.240000 ;
      RECT 0.000000 1670.790000 2368.360000 1671.690000 ;
      RECT 0.000000 1640.055000 2369.460000 1670.790000 ;
      RECT 1.100000 1639.155000 2369.460000 1640.055000 ;
      RECT 0.000000 1628.845000 2369.460000 1639.155000 ;
      RECT 0.000000 1627.945000 2368.360000 1628.845000 ;
      RECT 0.000000 1598.065000 2369.460000 1627.945000 ;
      RECT 1.100000 1597.165000 2369.460000 1598.065000 ;
      RECT 0.000000 1585.905000 2369.460000 1597.165000 ;
      RECT 0.000000 1585.005000 2368.360000 1585.905000 ;
      RECT 0.000000 1556.075000 2369.460000 1585.005000 ;
      RECT 1.100000 1555.175000 2369.460000 1556.075000 ;
      RECT 0.000000 1543.060000 2369.460000 1555.175000 ;
      RECT 0.000000 1542.160000 2368.360000 1543.060000 ;
      RECT 0.000000 1514.085000 2369.460000 1542.160000 ;
      RECT 1.100000 1513.185000 2369.460000 1514.085000 ;
      RECT 0.000000 1500.215000 2369.460000 1513.185000 ;
      RECT 0.000000 1499.315000 2368.360000 1500.215000 ;
      RECT 0.000000 1471.905000 2369.460000 1499.315000 ;
      RECT 1.100000 1471.005000 2369.460000 1471.905000 ;
      RECT 0.000000 1457.275000 2369.460000 1471.005000 ;
      RECT 0.000000 1456.375000 2368.360000 1457.275000 ;
      RECT 0.000000 1430.010000 2369.460000 1456.375000 ;
      RECT 1.100000 1429.110000 2369.460000 1430.010000 ;
      RECT 0.000000 1414.525000 2369.460000 1429.110000 ;
      RECT 0.000000 1413.625000 2368.360000 1414.525000 ;
      RECT 0.000000 1387.925000 2369.460000 1413.625000 ;
      RECT 1.100000 1387.025000 2369.460000 1387.925000 ;
      RECT 0.000000 1371.680000 2369.460000 1387.025000 ;
      RECT 0.000000 1370.780000 2368.360000 1371.680000 ;
      RECT 0.000000 1345.745000 2369.460000 1370.780000 ;
      RECT 1.100000 1344.845000 2369.460000 1345.745000 ;
      RECT 0.000000 1328.930000 2369.460000 1344.845000 ;
      RECT 0.000000 1328.030000 2368.360000 1328.930000 ;
      RECT 0.000000 1303.755000 2369.460000 1328.030000 ;
      RECT 1.100000 1302.855000 2369.460000 1303.755000 ;
      RECT 0.000000 1285.990000 2369.460000 1302.855000 ;
      RECT 0.000000 1285.090000 2368.360000 1285.990000 ;
      RECT 0.000000 1261.670000 2369.460000 1285.090000 ;
      RECT 1.100000 1260.770000 2369.460000 1261.670000 ;
      RECT 0.000000 1243.240000 2369.460000 1260.770000 ;
      RECT 0.000000 1242.340000 2368.360000 1243.240000 ;
      RECT 0.000000 1219.680000 2369.460000 1242.340000 ;
      RECT 1.100000 1218.780000 2369.460000 1219.680000 ;
      RECT 0.000000 1200.300000 2369.460000 1218.780000 ;
      RECT 0.000000 1199.400000 2368.360000 1200.300000 ;
      RECT 0.000000 1177.500000 2369.460000 1199.400000 ;
      RECT 1.100000 1176.600000 2369.460000 1177.500000 ;
      RECT 0.000000 1157.455000 2369.460000 1176.600000 ;
      RECT 0.000000 1156.555000 2368.360000 1157.455000 ;
      RECT 0.000000 1135.510000 2369.460000 1156.555000 ;
      RECT 1.100000 1134.610000 2369.460000 1135.510000 ;
      RECT 0.000000 1114.515000 2369.460000 1134.610000 ;
      RECT 0.000000 1113.615000 2368.360000 1114.515000 ;
      RECT 0.000000 1093.520000 2369.460000 1113.615000 ;
      RECT 1.100000 1092.620000 2369.460000 1093.520000 ;
      RECT 0.000000 1071.670000 2369.460000 1092.620000 ;
      RECT 0.000000 1070.770000 2368.360000 1071.670000 ;
      RECT 0.000000 1051.435000 2369.460000 1070.770000 ;
      RECT 1.100000 1050.535000 2369.460000 1051.435000 ;
      RECT 0.000000 1028.920000 2369.460000 1050.535000 ;
      RECT 0.000000 1028.020000 2368.360000 1028.920000 ;
      RECT 0.000000 1009.445000 2369.460000 1028.020000 ;
      RECT 1.100000 1008.545000 2369.460000 1009.445000 ;
      RECT 0.000000 985.980000 2369.460000 1008.545000 ;
      RECT 0.000000 985.080000 2368.360000 985.980000 ;
      RECT 0.000000 967.360000 2369.460000 985.080000 ;
      RECT 1.100000 966.460000 2369.460000 967.360000 ;
      RECT 0.000000 943.040000 2369.460000 966.460000 ;
      RECT 0.000000 942.140000 2368.360000 943.040000 ;
      RECT 0.000000 925.275000 2369.460000 942.140000 ;
      RECT 1.100000 924.375000 2369.460000 925.275000 ;
      RECT 0.000000 900.290000 2369.460000 924.375000 ;
      RECT 0.000000 899.390000 2368.360000 900.290000 ;
      RECT 0.000000 883.190000 2369.460000 899.390000 ;
      RECT 1.100000 882.290000 2369.460000 883.190000 ;
      RECT 0.000000 857.445000 2369.460000 882.290000 ;
      RECT 0.000000 856.545000 2368.360000 857.445000 ;
      RECT 0.000000 841.200000 2369.460000 856.545000 ;
      RECT 1.100000 840.300000 2369.460000 841.200000 ;
      RECT 0.000000 814.600000 2369.460000 840.300000 ;
      RECT 0.000000 813.700000 2368.360000 814.600000 ;
      RECT 0.000000 799.115000 2369.460000 813.700000 ;
      RECT 1.100000 798.215000 2369.460000 799.115000 ;
      RECT 0.000000 771.565000 2369.460000 798.215000 ;
      RECT 0.000000 770.665000 2368.360000 771.565000 ;
      RECT 0.000000 757.030000 2369.460000 770.665000 ;
      RECT 1.100000 756.130000 2369.460000 757.030000 ;
      RECT 0.000000 728.815000 2369.460000 756.130000 ;
      RECT 0.000000 727.915000 2368.360000 728.815000 ;
      RECT 0.000000 715.135000 2369.460000 727.915000 ;
      RECT 1.100000 714.235000 2369.460000 715.135000 ;
      RECT 0.000000 685.970000 2369.460000 714.235000 ;
      RECT 0.000000 685.070000 2368.360000 685.970000 ;
      RECT 0.000000 672.955000 2369.460000 685.070000 ;
      RECT 1.100000 672.055000 2369.460000 672.955000 ;
      RECT 0.000000 643.030000 2369.460000 672.055000 ;
      RECT 0.000000 642.130000 2368.360000 643.030000 ;
      RECT 0.000000 630.870000 2369.460000 642.130000 ;
      RECT 1.100000 629.970000 2369.460000 630.870000 ;
      RECT 0.000000 600.185000 2369.460000 629.970000 ;
      RECT 0.000000 599.285000 2368.360000 600.185000 ;
      RECT 0.000000 588.880000 2369.460000 599.285000 ;
      RECT 1.100000 587.980000 2369.460000 588.880000 ;
      RECT 0.000000 557.245000 2369.460000 587.980000 ;
      RECT 0.000000 556.345000 2368.360000 557.245000 ;
      RECT 0.000000 546.890000 2369.460000 556.345000 ;
      RECT 1.100000 545.990000 2369.460000 546.890000 ;
      RECT 0.000000 514.495000 2369.460000 545.990000 ;
      RECT 0.000000 513.595000 2368.360000 514.495000 ;
      RECT 0.000000 504.900000 2369.460000 513.595000 ;
      RECT 1.100000 504.000000 2369.460000 504.900000 ;
      RECT 0.000000 471.650000 2369.460000 504.000000 ;
      RECT 0.000000 470.750000 2368.360000 471.650000 ;
      RECT 0.000000 462.720000 2369.460000 470.750000 ;
      RECT 1.100000 461.820000 2369.460000 462.720000 ;
      RECT 0.000000 428.805000 2369.460000 461.820000 ;
      RECT 0.000000 427.905000 2368.360000 428.805000 ;
      RECT 0.000000 420.730000 2369.460000 427.905000 ;
      RECT 1.100000 419.830000 2369.460000 420.730000 ;
      RECT 0.000000 385.960000 2369.460000 419.830000 ;
      RECT 0.000000 385.060000 2368.360000 385.960000 ;
      RECT 0.000000 378.645000 2369.460000 385.060000 ;
      RECT 1.100000 377.745000 2369.460000 378.645000 ;
      RECT 0.000000 343.115000 2369.460000 377.745000 ;
      RECT 0.000000 342.215000 2368.360000 343.115000 ;
      RECT 0.000000 336.465000 2369.460000 342.215000 ;
      RECT 1.100000 335.565000 2369.460000 336.465000 ;
      RECT 0.000000 300.175000 2369.460000 335.565000 ;
      RECT 0.000000 299.275000 2368.360000 300.175000 ;
      RECT 0.000000 294.570000 2369.460000 299.275000 ;
      RECT 1.100000 293.670000 2369.460000 294.570000 ;
      RECT 0.000000 257.330000 2369.460000 293.670000 ;
      RECT 0.000000 256.430000 2368.360000 257.330000 ;
      RECT 0.000000 252.580000 2369.460000 256.430000 ;
      RECT 1.100000 251.680000 2369.460000 252.580000 ;
      RECT 0.000000 214.485000 2369.460000 251.680000 ;
      RECT 0.000000 213.585000 2368.360000 214.485000 ;
      RECT 0.000000 210.400000 2369.460000 213.585000 ;
      RECT 1.100000 209.500000 2369.460000 210.400000 ;
      RECT 0.000000 171.545000 2369.460000 209.500000 ;
      RECT 0.000000 170.645000 2368.360000 171.545000 ;
      RECT 0.000000 168.315000 2369.460000 170.645000 ;
      RECT 1.100000 167.415000 2369.460000 168.315000 ;
      RECT 0.000000 128.700000 2369.460000 167.415000 ;
      RECT 0.000000 127.800000 2368.360000 128.700000 ;
      RECT 0.000000 126.420000 2369.460000 127.800000 ;
      RECT 1.100000 125.520000 2369.460000 126.420000 ;
      RECT 0.000000 85.855000 2369.460000 125.520000 ;
      RECT 0.000000 84.955000 2368.360000 85.855000 ;
      RECT 0.000000 84.335000 2369.460000 84.955000 ;
      RECT 1.100000 83.435000 2369.460000 84.335000 ;
      RECT 0.000000 43.105000 2369.460000 83.435000 ;
      RECT 0.000000 42.250000 2368.360000 43.105000 ;
      RECT 1.100000 42.205000 2368.360000 42.250000 ;
      RECT 1.100000 41.350000 2369.460000 42.205000 ;
      RECT 0.000000 18.460000 2369.460000 41.350000 ;
      RECT 2356.080000 13.660000 2369.460000 18.460000 ;
      RECT 0.000000 13.660000 13.380000 18.460000 ;
      RECT 0.000000 12.660000 2369.460000 13.660000 ;
      RECT 2361.880000 7.860000 2369.460000 12.660000 ;
      RECT 0.000000 7.860000 7.580000 12.660000 ;
      RECT 0.000000 3.015000 2369.460000 7.860000 ;
      RECT 0.000000 2.255000 2368.360000 3.015000 ;
      RECT 1.100000 2.115000 2368.360000 2.255000 ;
      RECT 1.100000 1.355000 2369.460000 2.115000 ;
      RECT 0.000000 0.000000 2369.460000 1.355000 ;
    LAYER met4 ;
      RECT 0.000000 2281.700000 2369.460000 2290.240000 ;
      RECT 12.380000 2275.900000 2357.080000 2281.700000 ;
      RECT 2356.080000 13.660000 2357.080000 2275.900000 ;
      RECT 18.180000 13.660000 2351.280000 2275.900000 ;
      RECT 12.380000 13.660000 13.380000 2275.900000 ;
      RECT 2361.880000 7.860000 2369.460000 2281.700000 ;
      RECT 12.380000 7.860000 2357.080000 13.660000 ;
      RECT 0.000000 7.860000 7.580000 2281.700000 ;
      RECT 0.000000 0.000000 2369.460000 7.860000 ;
  END
END rest_top

END LIBRARY
