##
## LEF for PtnCells ;
## created by Innovus v20.10-p004_1 on Sat Dec 25 01:49:48 2021
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO rest_top
  CLASS BLOCK ;
  SIZE 2225.940000 BY 2895.100000 ;
  FOREIGN rest_top 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.430000 0.000000 4.570000 0.490000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.430000 0.000000 2.570000 0.485000 ;
    END
  END wb_rst_i
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.430000 0.000000 469.570000 0.490000 ;
    END
  END wbs_stb_i
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.930000 0.000000 158.070000 0.490000 ;
    END
  END wbs_cyc_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.930000 0.000000 474.070000 0.490000 ;
    END
  END wbs_we_i
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.930000 0.000000 465.070000 0.490000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.430000 0.000000 460.570000 0.490000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.930000 0.000000 456.070000 0.490000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.430000 0.000000 451.570000 0.490000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.430000 0.000000 302.570000 0.490000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.830000 0.000000 297.970000 0.490000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.330000 0.000000 293.470000 0.490000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.830000 0.000000 288.970000 0.490000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.330000 0.000000 284.470000 0.490000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.830000 0.000000 279.970000 0.490000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.330000 0.000000 275.470000 0.490000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.830000 0.000000 270.970000 0.490000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.230000 0.000000 266.370000 0.490000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.730000 0.000000 261.870000 0.490000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.230000 0.000000 257.370000 0.490000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.730000 0.000000 252.870000 0.490000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.230000 0.000000 248.370000 0.490000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.730000 0.000000 243.870000 0.490000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.130000 0.000000 239.270000 0.490000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.630000 0.000000 234.770000 0.490000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.130000 0.000000 230.270000 0.490000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.630000 0.000000 225.770000 0.490000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.130000 0.000000 221.270000 0.490000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.630000 0.000000 216.770000 0.490000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.130000 0.000000 212.270000 0.490000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.530000 0.000000 207.670000 0.490000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.030000 0.000000 203.170000 0.490000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.530000 0.000000 198.670000 0.490000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.030000 0.000000 194.170000 0.490000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.530000 0.000000 189.670000 0.490000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.030000 0.000000 185.170000 0.490000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.530000 0.000000 180.670000 0.490000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.930000 0.000000 176.070000 0.490000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.430000 0.000000 171.570000 0.490000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.930000 0.000000 167.070000 0.490000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.430000 0.000000 162.570000 0.490000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.430000 0.000000 153.570000 0.490000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.830000 0.000000 148.970000 0.490000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.330000 0.000000 144.470000 0.490000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.830000 0.000000 139.970000 0.490000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330000 0.000000 135.470000 0.490000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.830000 0.000000 130.970000 0.490000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.330000 0.000000 126.470000 0.490000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.830000 0.000000 121.970000 0.490000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.230000 0.000000 117.370000 0.490000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.730000 0.000000 112.870000 0.490000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.230000 0.000000 108.370000 0.490000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.730000 0.000000 103.870000 0.490000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.230000 0.000000 99.370000 0.490000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.730000 0.000000 94.870000 0.490000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.230000 0.000000 90.370000 0.490000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.630000 0.000000 85.770000 0.490000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.130000 0.000000 81.270000 0.490000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.630000 0.000000 76.770000 0.490000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.130000 0.000000 72.270000 0.490000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.630000 0.000000 67.770000 0.490000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.130000 0.000000 63.270000 0.490000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.530000 0.000000 58.670000 0.490000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.030000 0.000000 54.170000 0.490000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.530000 0.000000 49.670000 0.490000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.030000 0.000000 45.170000 0.490000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.530000 0.000000 40.670000 0.490000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.030000 0.000000 36.170000 0.490000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.530000 0.000000 31.670000 0.490000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.930000 0.000000 27.070000 0.490000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.430000 0.000000 22.570000 0.490000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.930000 0.000000 18.070000 0.490000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.430000 0.000000 13.570000 0.490000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_ack_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.930000 0.000000 9.070000 0.490000 ;
    END
  END wbs_ack_o
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.830000 0.000000 446.970000 0.490000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.330000 0.000000 442.470000 0.490000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.830000 0.000000 437.970000 0.490000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.330000 0.000000 433.470000 0.490000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.830000 0.000000 428.970000 0.490000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.330000 0.000000 424.470000 0.490000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.730000 0.000000 419.870000 0.490000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.230000 0.000000 415.370000 0.490000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.730000 0.000000 410.870000 0.490000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.230000 0.000000 406.370000 0.490000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.730000 0.000000 401.870000 0.490000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.230000 0.000000 397.370000 0.490000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.730000 0.000000 392.870000 0.490000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.130000 0.000000 388.270000 0.490000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.630000 0.000000 383.770000 0.490000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.130000 0.000000 379.270000 0.490000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.630000 0.000000 374.770000 0.490000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.130000 0.000000 370.270000 0.490000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.630000 0.000000 365.770000 0.490000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.130000 0.000000 361.270000 0.490000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.530000 0.000000 356.670000 0.490000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.030000 0.000000 352.170000 0.490000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.530000 0.000000 347.670000 0.490000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.030000 0.000000 343.170000 0.490000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.530000 0.000000 338.670000 0.490000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.030000 0.000000 334.170000 0.490000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.430000 0.000000 329.570000 0.490000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.930000 0.000000 325.070000 0.490000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.430000 0.000000 320.570000 0.490000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.930000 0.000000 316.070000 0.490000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.430000 0.000000 311.570000 0.490000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.930000 0.000000 307.070000 0.490000 ;
    END
  END wbs_dat_o[0]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1051.830000 0.000000 1051.970000 0.490000 ;
    END
  END la_data_in[127]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1047.330000 0.000000 1047.470000 0.490000 ;
    END
  END la_data_in[126]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1042.830000 0.000000 1042.970000 0.490000 ;
    END
  END la_data_in[125]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1038.330000 0.000000 1038.470000 0.490000 ;
    END
  END la_data_in[124]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1033.830000 0.000000 1033.970000 0.490000 ;
    END
  END la_data_in[123]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1029.330000 0.000000 1029.470000 0.490000 ;
    END
  END la_data_in[122]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.830000 0.000000 1024.970000 0.490000 ;
    END
  END la_data_in[121]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1020.230000 0.000000 1020.370000 0.490000 ;
    END
  END la_data_in[120]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1015.730000 0.000000 1015.870000 0.490000 ;
    END
  END la_data_in[119]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1011.230000 0.000000 1011.370000 0.490000 ;
    END
  END la_data_in[118]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1006.730000 0.000000 1006.870000 0.490000 ;
    END
  END la_data_in[117]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1002.230000 0.000000 1002.370000 0.490000 ;
    END
  END la_data_in[116]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 997.730000 0.000000 997.870000 0.490000 ;
    END
  END la_data_in[115]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 993.230000 0.000000 993.370000 0.490000 ;
    END
  END la_data_in[114]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 988.630000 0.000000 988.770000 0.490000 ;
    END
  END la_data_in[113]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 984.130000 0.000000 984.270000 0.490000 ;
    END
  END la_data_in[112]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 979.630000 0.000000 979.770000 0.490000 ;
    END
  END la_data_in[111]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 975.130000 0.000000 975.270000 0.490000 ;
    END
  END la_data_in[110]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 970.630000 0.000000 970.770000 0.490000 ;
    END
  END la_data_in[109]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 966.130000 0.000000 966.270000 0.490000 ;
    END
  END la_data_in[108]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 961.530000 0.000000 961.670000 0.490000 ;
    END
  END la_data_in[107]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 957.030000 0.000000 957.170000 0.490000 ;
    END
  END la_data_in[106]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 952.530000 0.000000 952.670000 0.490000 ;
    END
  END la_data_in[105]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.030000 0.000000 948.170000 0.490000 ;
    END
  END la_data_in[104]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 943.530000 0.000000 943.670000 0.490000 ;
    END
  END la_data_in[103]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 939.030000 0.000000 939.170000 0.490000 ;
    END
  END la_data_in[102]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 934.530000 0.000000 934.670000 0.490000 ;
    END
  END la_data_in[101]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 929.930000 0.000000 930.070000 0.490000 ;
    END
  END la_data_in[100]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 925.430000 0.000000 925.570000 0.490000 ;
    END
  END la_data_in[99]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 920.930000 0.000000 921.070000 0.490000 ;
    END
  END la_data_in[98]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 916.430000 0.000000 916.570000 0.490000 ;
    END
  END la_data_in[97]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.930000 0.000000 912.070000 0.490000 ;
    END
  END la_data_in[96]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.430000 0.000000 907.570000 0.490000 ;
    END
  END la_data_in[95]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 902.930000 0.000000 903.070000 0.490000 ;
    END
  END la_data_in[94]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.330000 0.000000 898.470000 0.490000 ;
    END
  END la_data_in[93]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 893.830000 0.000000 893.970000 0.490000 ;
    END
  END la_data_in[92]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.330000 0.000000 889.470000 0.490000 ;
    END
  END la_data_in[91]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 884.830000 0.000000 884.970000 0.490000 ;
    END
  END la_data_in[90]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 880.330000 0.000000 880.470000 0.490000 ;
    END
  END la_data_in[89]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.830000 0.000000 875.970000 0.490000 ;
    END
  END la_data_in[88]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.230000 0.000000 871.370000 0.490000 ;
    END
  END la_data_in[87]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 866.730000 0.000000 866.870000 0.490000 ;
    END
  END la_data_in[86]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 862.230000 0.000000 862.370000 0.490000 ;
    END
  END la_data_in[85]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 857.730000 0.000000 857.870000 0.490000 ;
    END
  END la_data_in[84]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.230000 0.000000 853.370000 0.490000 ;
    END
  END la_data_in[83]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 848.730000 0.000000 848.870000 0.490000 ;
    END
  END la_data_in[82]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 844.230000 0.000000 844.370000 0.490000 ;
    END
  END la_data_in[81]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 839.630000 0.000000 839.770000 0.490000 ;
    END
  END la_data_in[80]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.130000 0.000000 835.270000 0.490000 ;
    END
  END la_data_in[79]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.630000 0.000000 830.770000 0.490000 ;
    END
  END la_data_in[78]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 826.130000 0.000000 826.270000 0.490000 ;
    END
  END la_data_in[77]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.630000 0.000000 821.770000 0.490000 ;
    END
  END la_data_in[76]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.130000 0.000000 817.270000 0.490000 ;
    END
  END la_data_in[75]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 812.630000 0.000000 812.770000 0.490000 ;
    END
  END la_data_in[74]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 808.030000 0.000000 808.170000 0.490000 ;
    END
  END la_data_in[73]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 803.530000 0.000000 803.670000 0.490000 ;
    END
  END la_data_in[72]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 799.030000 0.000000 799.170000 0.490000 ;
    END
  END la_data_in[71]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.530000 0.000000 794.670000 0.490000 ;
    END
  END la_data_in[70]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 790.030000 0.000000 790.170000 0.490000 ;
    END
  END la_data_in[69]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.530000 0.000000 785.670000 0.490000 ;
    END
  END la_data_in[68]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 780.930000 0.000000 781.070000 0.490000 ;
    END
  END la_data_in[67]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.430000 0.000000 776.570000 0.490000 ;
    END
  END la_data_in[66]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.930000 0.000000 772.070000 0.490000 ;
    END
  END la_data_in[65]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.430000 0.000000 767.570000 0.490000 ;
    END
  END la_data_in[64]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 762.930000 0.000000 763.070000 0.490000 ;
    END
  END la_data_in[63]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.430000 0.000000 758.570000 0.490000 ;
    END
  END la_data_in[62]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.930000 0.000000 754.070000 0.490000 ;
    END
  END la_data_in[61]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.330000 0.000000 749.470000 0.490000 ;
    END
  END la_data_in[60]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 744.830000 0.000000 744.970000 0.490000 ;
    END
  END la_data_in[59]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.330000 0.000000 740.470000 0.490000 ;
    END
  END la_data_in[58]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.830000 0.000000 735.970000 0.490000 ;
    END
  END la_data_in[57]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.330000 0.000000 731.470000 0.490000 ;
    END
  END la_data_in[56]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 726.830000 0.000000 726.970000 0.490000 ;
    END
  END la_data_in[55]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.330000 0.000000 722.470000 0.490000 ;
    END
  END la_data_in[54]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.730000 0.000000 717.870000 0.490000 ;
    END
  END la_data_in[53]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.230000 0.000000 713.370000 0.490000 ;
    END
  END la_data_in[52]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.730000 0.000000 708.870000 0.490000 ;
    END
  END la_data_in[51]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.230000 0.000000 704.370000 0.490000 ;
    END
  END la_data_in[50]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.730000 0.000000 699.870000 0.490000 ;
    END
  END la_data_in[49]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.230000 0.000000 695.370000 0.490000 ;
    END
  END la_data_in[48]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.630000 0.000000 690.770000 0.490000 ;
    END
  END la_data_in[47]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.130000 0.000000 686.270000 0.490000 ;
    END
  END la_data_in[46]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 681.630000 0.000000 681.770000 0.490000 ;
    END
  END la_data_in[45]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 677.130000 0.000000 677.270000 0.490000 ;
    END
  END la_data_in[44]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.630000 0.000000 672.770000 0.490000 ;
    END
  END la_data_in[43]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.130000 0.000000 668.270000 0.490000 ;
    END
  END la_data_in[42]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.630000 0.000000 663.770000 0.490000 ;
    END
  END la_data_in[41]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 659.030000 0.000000 659.170000 0.490000 ;
    END
  END la_data_in[40]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 654.530000 0.000000 654.670000 0.490000 ;
    END
  END la_data_in[39]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.030000 0.000000 650.170000 0.490000 ;
    END
  END la_data_in[38]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.530000 0.000000 645.670000 0.490000 ;
    END
  END la_data_in[37]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.030000 0.000000 641.170000 0.490000 ;
    END
  END la_data_in[36]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 636.530000 0.000000 636.670000 0.490000 ;
    END
  END la_data_in[35]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.030000 0.000000 632.170000 0.490000 ;
    END
  END la_data_in[34]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.430000 0.000000 627.570000 0.490000 ;
    END
  END la_data_in[33]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.930000 0.000000 623.070000 0.490000 ;
    END
  END la_data_in[32]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.430000 0.000000 618.570000 0.490000 ;
    END
  END la_data_in[31]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 613.930000 0.000000 614.070000 0.490000 ;
    END
  END la_data_in[30]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.430000 0.000000 609.570000 0.490000 ;
    END
  END la_data_in[29]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.930000 0.000000 605.070000 0.490000 ;
    END
  END la_data_in[28]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 600.330000 0.000000 600.470000 0.490000 ;
    END
  END la_data_in[27]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.830000 0.000000 595.970000 0.490000 ;
    END
  END la_data_in[26]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.330000 0.000000 591.470000 0.490000 ;
    END
  END la_data_in[25]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.830000 0.000000 586.970000 0.490000 ;
    END
  END la_data_in[24]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.330000 0.000000 582.470000 0.490000 ;
    END
  END la_data_in[23]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.830000 0.000000 577.970000 0.490000 ;
    END
  END la_data_in[22]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.330000 0.000000 573.470000 0.490000 ;
    END
  END la_data_in[21]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 568.730000 0.000000 568.870000 0.490000 ;
    END
  END la_data_in[20]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.230000 0.000000 564.370000 0.490000 ;
    END
  END la_data_in[19]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.730000 0.000000 559.870000 0.490000 ;
    END
  END la_data_in[18]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.230000 0.000000 555.370000 0.490000 ;
    END
  END la_data_in[17]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.730000 0.000000 550.870000 0.490000 ;
    END
  END la_data_in[16]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.230000 0.000000 546.370000 0.490000 ;
    END
  END la_data_in[15]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.730000 0.000000 541.870000 0.490000 ;
    END
  END la_data_in[14]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.130000 0.000000 537.270000 0.490000 ;
    END
  END la_data_in[13]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.630000 0.000000 532.770000 0.490000 ;
    END
  END la_data_in[12]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.130000 0.000000 528.270000 0.490000 ;
    END
  END la_data_in[11]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.630000 0.000000 523.770000 0.490000 ;
    END
  END la_data_in[10]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.130000 0.000000 519.270000 0.490000 ;
    END
  END la_data_in[9]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.630000 0.000000 514.770000 0.490000 ;
    END
  END la_data_in[8]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.030000 0.000000 510.170000 0.490000 ;
    END
  END la_data_in[7]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.530000 0.000000 505.670000 0.490000 ;
    END
  END la_data_in[6]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.030000 0.000000 501.170000 0.490000 ;
    END
  END la_data_in[5]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.530000 0.000000 496.670000 0.490000 ;
    END
  END la_data_in[4]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.030000 0.000000 492.170000 0.490000 ;
    END
  END la_data_in[3]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.530000 0.000000 487.670000 0.490000 ;
    END
  END la_data_in[2]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.030000 0.000000 483.170000 0.490000 ;
    END
  END la_data_in[1]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.430000 0.000000 478.570000 0.490000 ;
    END
  END la_data_in[0]
  PIN la_data_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1629.830000 0.000000 1629.970000 0.490000 ;
    END
  END la_data_out[127]
  PIN la_data_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1625.330000 0.000000 1625.470000 0.490000 ;
    END
  END la_data_out[126]
  PIN la_data_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1620.730000 0.000000 1620.870000 0.490000 ;
    END
  END la_data_out[125]
  PIN la_data_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1616.230000 0.000000 1616.370000 0.490000 ;
    END
  END la_data_out[124]
  PIN la_data_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1611.730000 0.000000 1611.870000 0.490000 ;
    END
  END la_data_out[123]
  PIN la_data_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1607.230000 0.000000 1607.370000 0.490000 ;
    END
  END la_data_out[122]
  PIN la_data_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1602.730000 0.000000 1602.870000 0.490000 ;
    END
  END la_data_out[121]
  PIN la_data_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1598.230000 0.000000 1598.370000 0.490000 ;
    END
  END la_data_out[120]
  PIN la_data_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1593.630000 0.000000 1593.770000 0.490000 ;
    END
  END la_data_out[119]
  PIN la_data_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1589.130000 0.000000 1589.270000 0.490000 ;
    END
  END la_data_out[118]
  PIN la_data_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1584.630000 0.000000 1584.770000 0.490000 ;
    END
  END la_data_out[117]
  PIN la_data_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1580.130000 0.000000 1580.270000 0.490000 ;
    END
  END la_data_out[116]
  PIN la_data_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1575.630000 0.000000 1575.770000 0.490000 ;
    END
  END la_data_out[115]
  PIN la_data_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1571.130000 0.000000 1571.270000 0.490000 ;
    END
  END la_data_out[114]
  PIN la_data_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1566.630000 0.000000 1566.770000 0.490000 ;
    END
  END la_data_out[113]
  PIN la_data_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1562.030000 0.000000 1562.170000 0.490000 ;
    END
  END la_data_out[112]
  PIN la_data_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1557.530000 0.000000 1557.670000 0.490000 ;
    END
  END la_data_out[111]
  PIN la_data_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1553.030000 0.000000 1553.170000 0.490000 ;
    END
  END la_data_out[110]
  PIN la_data_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1548.530000 0.000000 1548.670000 0.490000 ;
    END
  END la_data_out[109]
  PIN la_data_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1544.030000 0.000000 1544.170000 0.490000 ;
    END
  END la_data_out[108]
  PIN la_data_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1539.530000 0.000000 1539.670000 0.490000 ;
    END
  END la_data_out[107]
  PIN la_data_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1535.030000 0.000000 1535.170000 0.490000 ;
    END
  END la_data_out[106]
  PIN la_data_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1530.430000 0.000000 1530.570000 0.490000 ;
    END
  END la_data_out[105]
  PIN la_data_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1525.930000 0.000000 1526.070000 0.490000 ;
    END
  END la_data_out[104]
  PIN la_data_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1521.430000 0.000000 1521.570000 0.490000 ;
    END
  END la_data_out[103]
  PIN la_data_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1516.930000 0.000000 1517.070000 0.490000 ;
    END
  END la_data_out[102]
  PIN la_data_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1512.430000 0.000000 1512.570000 0.490000 ;
    END
  END la_data_out[101]
  PIN la_data_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1507.930000 0.000000 1508.070000 0.490000 ;
    END
  END la_data_out[100]
  PIN la_data_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1503.330000 0.000000 1503.470000 0.490000 ;
    END
  END la_data_out[99]
  PIN la_data_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1498.830000 0.000000 1498.970000 0.490000 ;
    END
  END la_data_out[98]
  PIN la_data_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1494.330000 0.000000 1494.470000 0.490000 ;
    END
  END la_data_out[97]
  PIN la_data_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1489.830000 0.000000 1489.970000 0.490000 ;
    END
  END la_data_out[96]
  PIN la_data_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1485.330000 0.000000 1485.470000 0.490000 ;
    END
  END la_data_out[95]
  PIN la_data_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1480.830000 0.000000 1480.970000 0.490000 ;
    END
  END la_data_out[94]
  PIN la_data_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1476.330000 0.000000 1476.470000 0.490000 ;
    END
  END la_data_out[93]
  PIN la_data_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1471.730000 0.000000 1471.870000 0.490000 ;
    END
  END la_data_out[92]
  PIN la_data_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1467.230000 0.000000 1467.370000 0.490000 ;
    END
  END la_data_out[91]
  PIN la_data_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1462.730000 0.000000 1462.870000 0.490000 ;
    END
  END la_data_out[90]
  PIN la_data_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1458.230000 0.000000 1458.370000 0.490000 ;
    END
  END la_data_out[89]
  PIN la_data_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1453.730000 0.000000 1453.870000 0.490000 ;
    END
  END la_data_out[88]
  PIN la_data_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1449.230000 0.000000 1449.370000 0.490000 ;
    END
  END la_data_out[87]
  PIN la_data_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1444.730000 0.000000 1444.870000 0.490000 ;
    END
  END la_data_out[86]
  PIN la_data_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1440.130000 0.000000 1440.270000 0.490000 ;
    END
  END la_data_out[85]
  PIN la_data_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1435.630000 0.000000 1435.770000 0.490000 ;
    END
  END la_data_out[84]
  PIN la_data_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1431.130000 0.000000 1431.270000 0.490000 ;
    END
  END la_data_out[83]
  PIN la_data_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1426.630000 0.000000 1426.770000 0.490000 ;
    END
  END la_data_out[82]
  PIN la_data_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1422.130000 0.000000 1422.270000 0.490000 ;
    END
  END la_data_out[81]
  PIN la_data_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1417.630000 0.000000 1417.770000 0.490000 ;
    END
  END la_data_out[80]
  PIN la_data_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1413.030000 0.000000 1413.170000 0.490000 ;
    END
  END la_data_out[79]
  PIN la_data_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1408.530000 0.000000 1408.670000 0.490000 ;
    END
  END la_data_out[78]
  PIN la_data_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1404.030000 0.000000 1404.170000 0.490000 ;
    END
  END la_data_out[77]
  PIN la_data_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1399.530000 0.000000 1399.670000 0.490000 ;
    END
  END la_data_out[76]
  PIN la_data_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1395.030000 0.000000 1395.170000 0.490000 ;
    END
  END la_data_out[75]
  PIN la_data_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1390.530000 0.000000 1390.670000 0.490000 ;
    END
  END la_data_out[74]
  PIN la_data_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1386.030000 0.000000 1386.170000 0.490000 ;
    END
  END la_data_out[73]
  PIN la_data_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1381.430000 0.000000 1381.570000 0.490000 ;
    END
  END la_data_out[72]
  PIN la_data_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1376.930000 0.000000 1377.070000 0.490000 ;
    END
  END la_data_out[71]
  PIN la_data_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1372.430000 0.000000 1372.570000 0.490000 ;
    END
  END la_data_out[70]
  PIN la_data_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1367.930000 0.000000 1368.070000 0.490000 ;
    END
  END la_data_out[69]
  PIN la_data_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1363.430000 0.000000 1363.570000 0.490000 ;
    END
  END la_data_out[68]
  PIN la_data_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1358.930000 0.000000 1359.070000 0.490000 ;
    END
  END la_data_out[67]
  PIN la_data_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1354.430000 0.000000 1354.570000 0.490000 ;
    END
  END la_data_out[66]
  PIN la_data_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1349.830000 0.000000 1349.970000 0.490000 ;
    END
  END la_data_out[65]
  PIN la_data_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1345.330000 0.000000 1345.470000 0.490000 ;
    END
  END la_data_out[64]
  PIN la_data_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1340.830000 0.000000 1340.970000 0.490000 ;
    END
  END la_data_out[63]
  PIN la_data_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1336.330000 0.000000 1336.470000 0.490000 ;
    END
  END la_data_out[62]
  PIN la_data_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1331.830000 0.000000 1331.970000 0.490000 ;
    END
  END la_data_out[61]
  PIN la_data_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1327.330000 0.000000 1327.470000 0.490000 ;
    END
  END la_data_out[60]
  PIN la_data_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1322.730000 0.000000 1322.870000 0.490000 ;
    END
  END la_data_out[59]
  PIN la_data_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1318.230000 0.000000 1318.370000 0.490000 ;
    END
  END la_data_out[58]
  PIN la_data_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1313.730000 0.000000 1313.870000 0.490000 ;
    END
  END la_data_out[57]
  PIN la_data_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1309.230000 0.000000 1309.370000 0.490000 ;
    END
  END la_data_out[56]
  PIN la_data_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1304.730000 0.000000 1304.870000 0.490000 ;
    END
  END la_data_out[55]
  PIN la_data_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1300.230000 0.000000 1300.370000 0.490000 ;
    END
  END la_data_out[54]
  PIN la_data_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1295.730000 0.000000 1295.870000 0.490000 ;
    END
  END la_data_out[53]
  PIN la_data_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.130000 0.000000 1291.270000 0.490000 ;
    END
  END la_data_out[52]
  PIN la_data_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1286.630000 0.000000 1286.770000 0.490000 ;
    END
  END la_data_out[51]
  PIN la_data_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1282.130000 0.000000 1282.270000 0.490000 ;
    END
  END la_data_out[50]
  PIN la_data_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1277.630000 0.000000 1277.770000 0.490000 ;
    END
  END la_data_out[49]
  PIN la_data_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1273.130000 0.000000 1273.270000 0.490000 ;
    END
  END la_data_out[48]
  PIN la_data_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1268.630000 0.000000 1268.770000 0.490000 ;
    END
  END la_data_out[47]
  PIN la_data_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1264.130000 0.000000 1264.270000 0.490000 ;
    END
  END la_data_out[46]
  PIN la_data_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1259.530000 0.000000 1259.670000 0.490000 ;
    END
  END la_data_out[45]
  PIN la_data_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1255.030000 0.000000 1255.170000 0.490000 ;
    END
  END la_data_out[44]
  PIN la_data_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1250.530000 0.000000 1250.670000 0.490000 ;
    END
  END la_data_out[43]
  PIN la_data_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1246.030000 0.000000 1246.170000 0.490000 ;
    END
  END la_data_out[42]
  PIN la_data_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1241.530000 0.000000 1241.670000 0.490000 ;
    END
  END la_data_out[41]
  PIN la_data_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1237.030000 0.000000 1237.170000 0.490000 ;
    END
  END la_data_out[40]
  PIN la_data_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1232.430000 0.000000 1232.570000 0.490000 ;
    END
  END la_data_out[39]
  PIN la_data_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1227.930000 0.000000 1228.070000 0.490000 ;
    END
  END la_data_out[38]
  PIN la_data_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1223.430000 0.000000 1223.570000 0.490000 ;
    END
  END la_data_out[37]
  PIN la_data_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1218.930000 0.000000 1219.070000 0.490000 ;
    END
  END la_data_out[36]
  PIN la_data_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1214.430000 0.000000 1214.570000 0.490000 ;
    END
  END la_data_out[35]
  PIN la_data_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1209.930000 0.000000 1210.070000 0.490000 ;
    END
  END la_data_out[34]
  PIN la_data_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1205.430000 0.000000 1205.570000 0.490000 ;
    END
  END la_data_out[33]
  PIN la_data_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1200.830000 0.000000 1200.970000 0.490000 ;
    END
  END la_data_out[32]
  PIN la_data_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1196.330000 0.000000 1196.470000 0.490000 ;
    END
  END la_data_out[31]
  PIN la_data_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1191.830000 0.000000 1191.970000 0.490000 ;
    END
  END la_data_out[30]
  PIN la_data_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1187.330000 0.000000 1187.470000 0.490000 ;
    END
  END la_data_out[29]
  PIN la_data_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1182.830000 0.000000 1182.970000 0.490000 ;
    END
  END la_data_out[28]
  PIN la_data_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1178.330000 0.000000 1178.470000 0.490000 ;
    END
  END la_data_out[27]
  PIN la_data_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1173.830000 0.000000 1173.970000 0.490000 ;
    END
  END la_data_out[26]
  PIN la_data_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1169.230000 0.000000 1169.370000 0.490000 ;
    END
  END la_data_out[25]
  PIN la_data_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1164.730000 0.000000 1164.870000 0.490000 ;
    END
  END la_data_out[24]
  PIN la_data_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1160.230000 0.000000 1160.370000 0.490000 ;
    END
  END la_data_out[23]
  PIN la_data_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1155.730000 0.000000 1155.870000 0.490000 ;
    END
  END la_data_out[22]
  PIN la_data_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1151.230000 0.000000 1151.370000 0.490000 ;
    END
  END la_data_out[21]
  PIN la_data_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1146.730000 0.000000 1146.870000 0.490000 ;
    END
  END la_data_out[20]
  PIN la_data_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1142.130000 0.000000 1142.270000 0.490000 ;
    END
  END la_data_out[19]
  PIN la_data_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1137.630000 0.000000 1137.770000 0.490000 ;
    END
  END la_data_out[18]
  PIN la_data_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1133.130000 0.000000 1133.270000 0.490000 ;
    END
  END la_data_out[17]
  PIN la_data_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1128.630000 0.000000 1128.770000 0.490000 ;
    END
  END la_data_out[16]
  PIN la_data_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1124.130000 0.000000 1124.270000 0.490000 ;
    END
  END la_data_out[15]
  PIN la_data_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1119.630000 0.000000 1119.770000 0.490000 ;
    END
  END la_data_out[14]
  PIN la_data_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1115.130000 0.000000 1115.270000 0.490000 ;
    END
  END la_data_out[13]
  PIN la_data_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1110.530000 0.000000 1110.670000 0.490000 ;
    END
  END la_data_out[12]
  PIN la_data_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1106.030000 0.000000 1106.170000 0.490000 ;
    END
  END la_data_out[11]
  PIN la_data_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1101.530000 0.000000 1101.670000 0.490000 ;
    END
  END la_data_out[10]
  PIN la_data_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1097.030000 0.000000 1097.170000 0.490000 ;
    END
  END la_data_out[9]
  PIN la_data_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1092.530000 0.000000 1092.670000 0.490000 ;
    END
  END la_data_out[8]
  PIN la_data_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1088.030000 0.000000 1088.170000 0.490000 ;
    END
  END la_data_out[7]
  PIN la_data_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1083.530000 0.000000 1083.670000 0.490000 ;
    END
  END la_data_out[6]
  PIN la_data_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1078.930000 0.000000 1079.070000 0.490000 ;
    END
  END la_data_out[5]
  PIN la_data_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1074.430000 0.000000 1074.570000 0.490000 ;
    END
  END la_data_out[4]
  PIN la_data_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1069.930000 0.000000 1070.070000 0.490000 ;
    END
  END la_data_out[3]
  PIN la_data_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1065.430000 0.000000 1065.570000 0.490000 ;
    END
  END la_data_out[2]
  PIN la_data_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1060.930000 0.000000 1061.070000 0.490000 ;
    END
  END la_data_out[1]
  PIN la_data_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1056.430000 0.000000 1056.570000 0.490000 ;
    END
  END la_data_out[0]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2207.730000 0.000000 2207.870000 0.490000 ;
    END
  END la_oenb[127]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2203.230000 0.000000 2203.370000 0.490000 ;
    END
  END la_oenb[126]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2198.730000 0.000000 2198.870000 0.490000 ;
    END
  END la_oenb[125]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2194.130000 0.000000 2194.270000 0.490000 ;
    END
  END la_oenb[124]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2189.630000 0.000000 2189.770000 0.490000 ;
    END
  END la_oenb[123]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2185.130000 0.000000 2185.270000 0.490000 ;
    END
  END la_oenb[122]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2180.630000 0.000000 2180.770000 0.490000 ;
    END
  END la_oenb[121]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2176.130000 0.000000 2176.270000 0.490000 ;
    END
  END la_oenb[120]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2171.630000 0.000000 2171.770000 0.490000 ;
    END
  END la_oenb[119]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2167.130000 0.000000 2167.270000 0.490000 ;
    END
  END la_oenb[118]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2162.530000 0.000000 2162.670000 0.490000 ;
    END
  END la_oenb[117]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2158.030000 0.000000 2158.170000 0.490000 ;
    END
  END la_oenb[116]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2153.530000 0.000000 2153.670000 0.490000 ;
    END
  END la_oenb[115]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2149.030000 0.000000 2149.170000 0.490000 ;
    END
  END la_oenb[114]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2144.530000 0.000000 2144.670000 0.490000 ;
    END
  END la_oenb[113]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2140.030000 0.000000 2140.170000 0.490000 ;
    END
  END la_oenb[112]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2135.430000 0.000000 2135.570000 0.490000 ;
    END
  END la_oenb[111]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2130.930000 0.000000 2131.070000 0.490000 ;
    END
  END la_oenb[110]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2126.430000 0.000000 2126.570000 0.490000 ;
    END
  END la_oenb[109]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2121.930000 0.000000 2122.070000 0.490000 ;
    END
  END la_oenb[108]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2117.430000 0.000000 2117.570000 0.490000 ;
    END
  END la_oenb[107]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2112.930000 0.000000 2113.070000 0.490000 ;
    END
  END la_oenb[106]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2108.430000 0.000000 2108.570000 0.490000 ;
    END
  END la_oenb[105]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2103.830000 0.000000 2103.970000 0.490000 ;
    END
  END la_oenb[104]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2099.330000 0.000000 2099.470000 0.490000 ;
    END
  END la_oenb[103]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2094.830000 0.000000 2094.970000 0.490000 ;
    END
  END la_oenb[102]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2090.330000 0.000000 2090.470000 0.490000 ;
    END
  END la_oenb[101]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2085.830000 0.000000 2085.970000 0.490000 ;
    END
  END la_oenb[100]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2081.330000 0.000000 2081.470000 0.490000 ;
    END
  END la_oenb[99]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2076.830000 0.000000 2076.970000 0.490000 ;
    END
  END la_oenb[98]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2072.230000 0.000000 2072.370000 0.490000 ;
    END
  END la_oenb[97]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2067.730000 0.000000 2067.870000 0.490000 ;
    END
  END la_oenb[96]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2063.230000 0.000000 2063.370000 0.490000 ;
    END
  END la_oenb[95]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2058.730000 0.000000 2058.870000 0.490000 ;
    END
  END la_oenb[94]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2054.230000 0.000000 2054.370000 0.490000 ;
    END
  END la_oenb[93]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2049.730000 0.000000 2049.870000 0.490000 ;
    END
  END la_oenb[92]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2045.130000 0.000000 2045.270000 0.490000 ;
    END
  END la_oenb[91]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2040.630000 0.000000 2040.770000 0.490000 ;
    END
  END la_oenb[90]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2036.130000 0.000000 2036.270000 0.490000 ;
    END
  END la_oenb[89]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2031.630000 0.000000 2031.770000 0.490000 ;
    END
  END la_oenb[88]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2027.130000 0.000000 2027.270000 0.490000 ;
    END
  END la_oenb[87]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2022.630000 0.000000 2022.770000 0.490000 ;
    END
  END la_oenb[86]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2018.130000 0.000000 2018.270000 0.490000 ;
    END
  END la_oenb[85]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2013.530000 0.000000 2013.670000 0.490000 ;
    END
  END la_oenb[84]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2009.030000 0.000000 2009.170000 0.490000 ;
    END
  END la_oenb[83]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2004.530000 0.000000 2004.670000 0.490000 ;
    END
  END la_oenb[82]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2000.030000 0.000000 2000.170000 0.490000 ;
    END
  END la_oenb[81]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1995.530000 0.000000 1995.670000 0.490000 ;
    END
  END la_oenb[80]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1991.030000 0.000000 1991.170000 0.490000 ;
    END
  END la_oenb[79]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1986.530000 0.000000 1986.670000 0.490000 ;
    END
  END la_oenb[78]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1981.930000 0.000000 1982.070000 0.490000 ;
    END
  END la_oenb[77]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1977.430000 0.000000 1977.570000 0.490000 ;
    END
  END la_oenb[76]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1972.930000 0.000000 1973.070000 0.490000 ;
    END
  END la_oenb[75]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1968.430000 0.000000 1968.570000 0.490000 ;
    END
  END la_oenb[74]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1963.930000 0.000000 1964.070000 0.490000 ;
    END
  END la_oenb[73]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1959.430000 0.000000 1959.570000 0.490000 ;
    END
  END la_oenb[72]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1954.830000 0.000000 1954.970000 0.490000 ;
    END
  END la_oenb[71]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1950.330000 0.000000 1950.470000 0.490000 ;
    END
  END la_oenb[70]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1945.830000 0.000000 1945.970000 0.490000 ;
    END
  END la_oenb[69]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1941.330000 0.000000 1941.470000 0.490000 ;
    END
  END la_oenb[68]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1936.830000 0.000000 1936.970000 0.490000 ;
    END
  END la_oenb[67]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1932.330000 0.000000 1932.470000 0.490000 ;
    END
  END la_oenb[66]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1927.830000 0.000000 1927.970000 0.490000 ;
    END
  END la_oenb[65]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1923.230000 0.000000 1923.370000 0.490000 ;
    END
  END la_oenb[64]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1918.730000 0.000000 1918.870000 0.490000 ;
    END
  END la_oenb[63]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1914.230000 0.000000 1914.370000 0.490000 ;
    END
  END la_oenb[62]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1909.730000 0.000000 1909.870000 0.490000 ;
    END
  END la_oenb[61]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.230000 0.000000 1905.370000 0.490000 ;
    END
  END la_oenb[60]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1900.730000 0.000000 1900.870000 0.490000 ;
    END
  END la_oenb[59]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1896.230000 0.000000 1896.370000 0.490000 ;
    END
  END la_oenb[58]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1891.630000 0.000000 1891.770000 0.490000 ;
    END
  END la_oenb[57]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1887.130000 0.000000 1887.270000 0.490000 ;
    END
  END la_oenb[56]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1882.630000 0.000000 1882.770000 0.490000 ;
    END
  END la_oenb[55]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1878.130000 0.000000 1878.270000 0.490000 ;
    END
  END la_oenb[54]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1873.630000 0.000000 1873.770000 0.490000 ;
    END
  END la_oenb[53]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1869.130000 0.000000 1869.270000 0.490000 ;
    END
  END la_oenb[52]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1864.530000 0.000000 1864.670000 0.490000 ;
    END
  END la_oenb[51]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1860.030000 0.000000 1860.170000 0.490000 ;
    END
  END la_oenb[50]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1855.530000 0.000000 1855.670000 0.490000 ;
    END
  END la_oenb[49]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1851.030000 0.000000 1851.170000 0.490000 ;
    END
  END la_oenb[48]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1846.530000 0.000000 1846.670000 0.490000 ;
    END
  END la_oenb[47]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1842.030000 0.000000 1842.170000 0.490000 ;
    END
  END la_oenb[46]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1837.530000 0.000000 1837.670000 0.490000 ;
    END
  END la_oenb[45]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1832.930000 0.000000 1833.070000 0.490000 ;
    END
  END la_oenb[44]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1828.430000 0.000000 1828.570000 0.490000 ;
    END
  END la_oenb[43]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1823.930000 0.000000 1824.070000 0.490000 ;
    END
  END la_oenb[42]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1819.430000 0.000000 1819.570000 0.490000 ;
    END
  END la_oenb[41]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1814.930000 0.000000 1815.070000 0.490000 ;
    END
  END la_oenb[40]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1810.430000 0.000000 1810.570000 0.490000 ;
    END
  END la_oenb[39]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1805.930000 0.000000 1806.070000 0.490000 ;
    END
  END la_oenb[38]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1801.330000 0.000000 1801.470000 0.490000 ;
    END
  END la_oenb[37]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1796.830000 0.000000 1796.970000 0.490000 ;
    END
  END la_oenb[36]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1792.330000 0.000000 1792.470000 0.490000 ;
    END
  END la_oenb[35]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1787.830000 0.000000 1787.970000 0.490000 ;
    END
  END la_oenb[34]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1783.330000 0.000000 1783.470000 0.490000 ;
    END
  END la_oenb[33]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1778.830000 0.000000 1778.970000 0.490000 ;
    END
  END la_oenb[32]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1774.230000 0.000000 1774.370000 0.490000 ;
    END
  END la_oenb[31]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1769.730000 0.000000 1769.870000 0.490000 ;
    END
  END la_oenb[30]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1765.230000 0.000000 1765.370000 0.490000 ;
    END
  END la_oenb[29]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1760.730000 0.000000 1760.870000 0.490000 ;
    END
  END la_oenb[28]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1756.230000 0.000000 1756.370000 0.490000 ;
    END
  END la_oenb[27]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1751.730000 0.000000 1751.870000 0.490000 ;
    END
  END la_oenb[26]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1747.230000 0.000000 1747.370000 0.490000 ;
    END
  END la_oenb[25]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1742.630000 0.000000 1742.770000 0.490000 ;
    END
  END la_oenb[24]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1738.130000 0.000000 1738.270000 0.490000 ;
    END
  END la_oenb[23]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1733.630000 0.000000 1733.770000 0.490000 ;
    END
  END la_oenb[22]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1729.130000 0.000000 1729.270000 0.490000 ;
    END
  END la_oenb[21]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1724.630000 0.000000 1724.770000 0.490000 ;
    END
  END la_oenb[20]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1720.130000 0.000000 1720.270000 0.490000 ;
    END
  END la_oenb[19]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1715.630000 0.000000 1715.770000 0.490000 ;
    END
  END la_oenb[18]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1711.030000 0.000000 1711.170000 0.490000 ;
    END
  END la_oenb[17]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1706.530000 0.000000 1706.670000 0.490000 ;
    END
  END la_oenb[16]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1702.030000 0.000000 1702.170000 0.490000 ;
    END
  END la_oenb[15]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1697.530000 0.000000 1697.670000 0.490000 ;
    END
  END la_oenb[14]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1693.030000 0.000000 1693.170000 0.490000 ;
    END
  END la_oenb[13]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1688.530000 0.000000 1688.670000 0.490000 ;
    END
  END la_oenb[12]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1683.930000 0.000000 1684.070000 0.490000 ;
    END
  END la_oenb[11]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1679.430000 0.000000 1679.570000 0.490000 ;
    END
  END la_oenb[10]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1674.930000 0.000000 1675.070000 0.490000 ;
    END
  END la_oenb[9]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1670.430000 0.000000 1670.570000 0.490000 ;
    END
  END la_oenb[8]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1665.930000 0.000000 1666.070000 0.490000 ;
    END
  END la_oenb[7]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1661.430000 0.000000 1661.570000 0.490000 ;
    END
  END la_oenb[6]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1656.930000 0.000000 1657.070000 0.490000 ;
    END
  END la_oenb[5]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1652.330000 0.000000 1652.470000 0.490000 ;
    END
  END la_oenb[4]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1647.830000 0.000000 1647.970000 0.490000 ;
    END
  END la_oenb[3]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1643.330000 0.000000 1643.470000 0.490000 ;
    END
  END la_oenb[2]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1638.830000 0.000000 1638.970000 0.490000 ;
    END
  END la_oenb[1]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1634.330000 0.000000 1634.470000 0.490000 ;
    END
  END la_oenb[0]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 108.730000 0.800000 109.030000 ;
    END
  END io_in[37]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 272.095000 0.800000 272.395000 ;
    END
  END io_in[36]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 435.460000 0.800000 435.760000 ;
    END
  END io_in[35]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 653.315000 0.800000 653.615000 ;
    END
  END io_in[34]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 871.070000 0.800000 871.370000 ;
    END
  END io_in[33]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1088.925000 0.800000 1089.225000 ;
    END
  END io_in[32]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1306.780000 0.800000 1307.080000 ;
    END
  END io_in[31]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1524.535000 0.800000 1524.835000 ;
    END
  END io_in[30]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1742.390000 0.800000 1742.690000 ;
    END
  END io_in[29]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1960.240000 0.800000 1960.540000 ;
    END
  END io_in[28]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2178.000000 0.800000 2178.300000 ;
    END
  END io_in[27]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2395.850000 0.800000 2396.150000 ;
    END
  END io_in[26]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2613.705000 0.800000 2614.005000 ;
    END
  END io_in[25]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2831.460000 0.800000 2831.760000 ;
    END
  END io_in[24]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.030000 2894.610000 127.170000 2895.100000 ;
    END
  END io_in[23]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.430000 2894.610000 381.570000 2895.100000 ;
    END
  END io_in[22]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 635.830000 2894.610000 635.970000 2895.100000 ;
    END
  END io_in[21]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 890.230000 2894.610000 890.370000 2895.100000 ;
    END
  END io_in[20]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1144.630000 2894.610000 1144.770000 2895.100000 ;
    END
  END io_in[19]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1399.030000 2894.610000 1399.170000 2895.100000 ;
    END
  END io_in[18]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1653.430000 2894.610000 1653.570000 2895.100000 ;
    END
  END io_in[17]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1907.830000 2894.610000 1907.970000 2895.100000 ;
    END
  END io_in[16]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2162.230000 2894.610000 2162.370000 2895.100000 ;
    END
  END io_in[15]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 2775.015000 2225.940000 2775.315000 ;
    END
  END io_in[14]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 2552.945000 2225.940000 2553.245000 ;
    END
  END io_in[13]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 2330.975000 2225.940000 2331.275000 ;
    END
  END io_in[12]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 2108.910000 2225.940000 2109.210000 ;
    END
  END io_in[11]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 1886.940000 2225.940000 1887.240000 ;
    END
  END io_in[10]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 1664.870000 2225.940000 1665.170000 ;
    END
  END io_in[9]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 1442.900000 2225.940000 1443.200000 ;
    END
  END io_in[8]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 1220.830000 2225.940000 1221.130000 ;
    END
  END io_in[7]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 998.860000 2225.940000 999.160000 ;
    END
  END io_in[6]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 832.360000 2225.940000 832.660000 ;
    END
  END io_in[5]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 665.860000 2225.940000 666.160000 ;
    END
  END io_in[4]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 499.355000 2225.940000 499.655000 ;
    END
  END io_in[3]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 332.855000 2225.940000 333.155000 ;
    END
  END io_in[2]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 166.350000 2225.940000 166.650000 ;
    END
  END io_in[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 2.300000 2225.940000 2.600000 ;
    END
  END io_in[0]
  PIN io_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 54.240000 0.800000 54.540000 ;
    END
  END io_out[37]
  PIN io_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 217.605000 0.800000 217.905000 ;
    END
  END io_out[36]
  PIN io_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 380.970000 0.800000 381.270000 ;
    END
  END io_out[35]
  PIN io_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 598.825000 0.800000 599.125000 ;
    END
  END io_out[34]
  PIN io_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 816.680000 0.800000 816.980000 ;
    END
  END io_out[33]
  PIN io_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1034.435000 0.800000 1034.735000 ;
    END
  END io_out[32]
  PIN io_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1252.290000 0.800000 1252.590000 ;
    END
  END io_out[31]
  PIN io_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1470.145000 0.800000 1470.445000 ;
    END
  END io_out[30]
  PIN io_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1687.900000 0.800000 1688.200000 ;
    END
  END io_out[29]
  PIN io_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1905.755000 0.800000 1906.055000 ;
    END
  END io_out[28]
  PIN io_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2123.610000 0.800000 2123.910000 ;
    END
  END io_out[27]
  PIN io_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2341.365000 0.800000 2341.665000 ;
    END
  END io_out[26]
  PIN io_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2559.220000 0.800000 2559.520000 ;
    END
  END io_out[25]
  PIN io_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2777.070000 0.800000 2777.370000 ;
    END
  END io_out[24]
  PIN io_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.530000 2894.610000 63.670000 2895.100000 ;
    END
  END io_out[23]
  PIN io_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.830000 2894.610000 317.970000 2895.100000 ;
    END
  END io_out[22]
  PIN io_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.230000 2894.610000 572.370000 2895.100000 ;
    END
  END io_out[21]
  PIN io_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 826.630000 2894.610000 826.770000 2895.100000 ;
    END
  END io_out[20]
  PIN io_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1081.030000 2894.610000 1081.170000 2895.100000 ;
    END
  END io_out[19]
  PIN io_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1335.430000 2894.610000 1335.570000 2895.100000 ;
    END
  END io_out[18]
  PIN io_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1589.830000 2894.610000 1589.970000 2895.100000 ;
    END
  END io_out[17]
  PIN io_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1844.230000 2894.610000 1844.370000 2895.100000 ;
    END
  END io_out[16]
  PIN io_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2098.630000 2894.610000 2098.770000 2895.100000 ;
    END
  END io_out[15]
  PIN io_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 2830.480000 2225.940000 2830.780000 ;
    END
  END io_out[14]
  PIN io_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 2608.415000 2225.940000 2608.715000 ;
    END
  END io_out[13]
  PIN io_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 2386.445000 2225.940000 2386.745000 ;
    END
  END io_out[12]
  PIN io_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 2164.475000 2225.940000 2164.775000 ;
    END
  END io_out[11]
  PIN io_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 1942.405000 2225.940000 1942.705000 ;
    END
  END io_out[10]
  PIN io_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 1720.435000 2225.940000 1720.735000 ;
    END
  END io_out[9]
  PIN io_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 1498.370000 2225.940000 1498.670000 ;
    END
  END io_out[8]
  PIN io_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 1276.400000 2225.940000 1276.700000 ;
    END
  END io_out[7]
  PIN io_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 1054.330000 2225.940000 1054.630000 ;
    END
  END io_out[6]
  PIN io_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 887.830000 2225.940000 888.130000 ;
    END
  END io_out[5]
  PIN io_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 721.325000 2225.940000 721.625000 ;
    END
  END io_out[4]
  PIN io_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 554.825000 2225.940000 555.125000 ;
    END
  END io_out[3]
  PIN io_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 388.320000 2225.940000 388.620000 ;
    END
  END io_out[2]
  PIN io_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 221.820000 2225.940000 222.120000 ;
    END
  END io_out[1]
  PIN io_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 55.320000 2225.940000 55.620000 ;
    END
  END io_out[0]
  PIN io_oeb[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1.125000 0.800000 1.425000 ;
    END
  END io_oeb[37]
  PIN io_oeb[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 163.215000 0.800000 163.515000 ;
    END
  END io_oeb[36]
  PIN io_oeb[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 326.580000 0.800000 326.880000 ;
    END
  END io_oeb[35]
  PIN io_oeb[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 544.340000 0.800000 544.640000 ;
    END
  END io_oeb[34]
  PIN io_oeb[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 762.190000 0.800000 762.490000 ;
    END
  END io_oeb[33]
  PIN io_oeb[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 980.045000 0.800000 980.345000 ;
    END
  END io_oeb[32]
  PIN io_oeb[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1197.800000 0.800000 1198.100000 ;
    END
  END io_oeb[31]
  PIN io_oeb[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1415.655000 0.800000 1415.955000 ;
    END
  END io_oeb[30]
  PIN io_oeb[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1633.510000 0.800000 1633.810000 ;
    END
  END io_oeb[29]
  PIN io_oeb[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1851.265000 0.800000 1851.565000 ;
    END
  END io_oeb[28]
  PIN io_oeb[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2069.120000 0.800000 2069.420000 ;
    END
  END io_oeb[27]
  PIN io_oeb[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2286.975000 0.800000 2287.275000 ;
    END
  END io_oeb[26]
  PIN io_oeb[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2504.730000 0.800000 2505.030000 ;
    END
  END io_oeb[25]
  PIN io_oeb[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2722.585000 0.800000 2722.885000 ;
    END
  END io_oeb[24]
  PIN io_oeb[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.230000 2894.615000 4.370000 2895.100000 ;
    END
  END io_oeb[23]
  PIN io_oeb[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.230000 2894.610000 254.370000 2895.100000 ;
    END
  END io_oeb[22]
  PIN io_oeb[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.630000 2894.610000 508.770000 2895.100000 ;
    END
  END io_oeb[21]
  PIN io_oeb[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.030000 2894.610000 763.170000 2895.100000 ;
    END
  END io_oeb[20]
  PIN io_oeb[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1017.430000 2894.610000 1017.570000 2895.100000 ;
    END
  END io_oeb[19]
  PIN io_oeb[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1271.830000 2894.610000 1271.970000 2895.100000 ;
    END
  END io_oeb[18]
  PIN io_oeb[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1526.230000 2894.610000 1526.370000 2895.100000 ;
    END
  END io_oeb[17]
  PIN io_oeb[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1780.630000 2894.610000 1780.770000 2895.100000 ;
    END
  END io_oeb[16]
  PIN io_oeb[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2035.030000 2894.610000 2035.170000 2895.100000 ;
    END
  END io_oeb[15]
  PIN io_oeb[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 2883.695000 2225.940000 2883.995000 ;
    END
  END io_oeb[14]
  PIN io_oeb[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 2663.980000 2225.940000 2664.280000 ;
    END
  END io_oeb[13]
  PIN io_oeb[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 2441.910000 2225.940000 2442.210000 ;
    END
  END io_oeb[12]
  PIN io_oeb[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 2219.940000 2225.940000 2220.240000 ;
    END
  END io_oeb[11]
  PIN io_oeb[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 1997.875000 2225.940000 1998.175000 ;
    END
  END io_oeb[10]
  PIN io_oeb[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 1775.905000 2225.940000 1776.205000 ;
    END
  END io_oeb[9]
  PIN io_oeb[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 1553.935000 2225.940000 1554.235000 ;
    END
  END io_oeb[8]
  PIN io_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 1331.865000 2225.940000 1332.165000 ;
    END
  END io_oeb[7]
  PIN io_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 1109.895000 2225.940000 1110.195000 ;
    END
  END io_oeb[6]
  PIN io_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 943.395000 2225.940000 943.695000 ;
    END
  END io_oeb[5]
  PIN io_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 776.890000 2225.940000 777.190000 ;
    END
  END io_oeb[4]
  PIN io_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 610.290000 2225.940000 610.590000 ;
    END
  END io_oeb[3]
  PIN io_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 443.790000 2225.940000 444.090000 ;
    END
  END io_oeb[2]
  PIN io_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 277.290000 2225.940000 277.590000 ;
    END
  END io_oeb[1]
  PIN io_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 110.785000 2225.940000 111.085000 ;
    END
  END io_oeb[0]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 489.950000 0.800000 490.250000 ;
    END
  END analog_io[28]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 707.705000 0.800000 708.005000 ;
    END
  END analog_io[27]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 925.560000 0.800000 925.860000 ;
    END
  END analog_io[26]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1143.410000 0.800000 1143.710000 ;
    END
  END analog_io[25]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1361.170000 0.800000 1361.470000 ;
    END
  END analog_io[24]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1579.020000 0.800000 1579.320000 ;
    END
  END analog_io[23]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1796.875000 0.800000 1797.175000 ;
    END
  END analog_io[22]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2014.630000 0.800000 2014.930000 ;
    END
  END analog_io[21]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2232.485000 0.800000 2232.785000 ;
    END
  END analog_io[20]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2450.340000 0.800000 2450.640000 ;
    END
  END analog_io[19]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2668.095000 0.800000 2668.395000 ;
    END
  END analog_io[18]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2883.110000 0.800000 2883.410000 ;
    END
  END analog_io[17]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.630000 2894.610000 190.770000 2895.100000 ;
    END
  END analog_io[16]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.030000 2894.610000 445.170000 2895.100000 ;
    END
  END analog_io[15]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.430000 2894.610000 699.570000 2895.100000 ;
    END
  END analog_io[14]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.830000 2894.610000 953.970000 2895.100000 ;
    END
  END analog_io[13]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1208.230000 2894.610000 1208.370000 2895.100000 ;
    END
  END analog_io[12]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1462.630000 2894.610000 1462.770000 2895.100000 ;
    END
  END analog_io[11]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1717.030000 2894.610000 1717.170000 2895.100000 ;
    END
  END analog_io[10]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1971.430000 2894.610000 1971.570000 2895.100000 ;
    END
  END analog_io[9]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2222.330000 2894.615000 2222.470000 2895.100000 ;
    END
  END analog_io[8]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 2719.450000 2225.940000 2719.750000 ;
    END
  END analog_io[7]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 2497.480000 2225.940000 2497.780000 ;
    END
  END analog_io[6]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 2275.410000 2225.940000 2275.710000 ;
    END
  END analog_io[5]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 2053.440000 2225.940000 2053.740000 ;
    END
  END analog_io[4]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 1831.370000 2225.940000 1831.670000 ;
    END
  END analog_io[3]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 1609.400000 2225.940000 1609.700000 ;
    END
  END analog_io[2]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 1387.430000 2225.940000 1387.730000 ;
    END
  END analog_io[1]
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2225.140000 1165.365000 2225.940000 1165.665000 ;
    END
  END analog_io[0]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2212.230000 0.000000 2212.370000 0.490000 ;
    END
  END user_clock2
  PIN user_irq[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2224.230000 0.000000 2224.370000 0.485000 ;
    END
  END user_irq[2]
  PIN user_irq[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2221.230000 0.000000 2221.370000 0.490000 ;
    END
  END user_irq[1]
  PIN user_irq[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2216.730000 0.000000 2216.870000 0.490000 ;
    END
  END user_irq[0]
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 7.980000 8.260000 2217.960000 12.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.980000 2881.140000 2217.960000 2885.140000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2213.960000 8.260000 2217.960000 2885.140000 ;
    END
    PORT
      LAYER met4 ;
        RECT 7.980000 8.260000 11.980000 2885.140000 ;
    END

# P/G pin shape extracted from block 'tcam_32x28'
    PORT
      LAYER met4 ;
        RECT 1109.555000 2373.635000 1111.295000 2768.415000 ;
      LAYER met3 ;
        RECT 1109.555000 2766.675000 1586.615000 2768.415000 ;
      LAYER met3 ;
        RECT 1109.555000 2373.635000 1586.615000 2375.375000 ;
      LAYER met4 ;
        RECT 1584.875000 2373.635000 1586.615000 2768.415000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1671.695000 2373.730000 1673.435000 2768.510000 ;
      LAYER met3 ;
        RECT 1671.695000 2766.770000 2148.755000 2768.510000 ;
      LAYER met3 ;
        RECT 1671.695000 2373.730000 2148.755000 2375.470000 ;
      LAYER met4 ;
        RECT 2147.015000 2373.730000 2148.755000 2768.510000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1083.485000 2334.200000 1085.485000 2804.040000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2173.025000 2334.200000 2175.025000 2804.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1083.485000 2802.040000 2175.025000 2804.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1083.485000 2334.200000 2175.025000 2336.200000 ;
    END
# end of P/G pin shape extracted from block 'tcam_32x28'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1556.385000 350.985000 1558.125000 745.765000 ;
      LAYER met3 ;
        RECT 1081.065000 350.985000 1558.125000 352.725000 ;
      LAYER met3 ;
        RECT 1081.065000 744.025000 1558.125000 745.765000 ;
      LAYER met4 ;
        RECT 1081.065000 350.985000 1082.805000 745.765000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1556.385000 848.485000 1558.125000 1243.265000 ;
      LAYER met3 ;
        RECT 1081.065000 848.485000 1558.125000 850.225000 ;
      LAYER met3 ;
        RECT 1081.065000 1241.525000 1558.125000 1243.265000 ;
      LAYER met4 ;
        RECT 1081.065000 848.485000 1082.805000 1243.265000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1556.385000 1843.485000 1558.125000 2238.265000 ;
      LAYER met3 ;
        RECT 1081.065000 1843.485000 1558.125000 1845.225000 ;
      LAYER met3 ;
        RECT 1081.065000 2236.525000 1558.125000 2238.265000 ;
      LAYER met4 ;
        RECT 1081.065000 1843.485000 1082.805000 2238.265000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1556.385000 1345.985000 1558.125000 1740.765000 ;
      LAYER met3 ;
        RECT 1081.065000 1345.985000 1558.125000 1347.725000 ;
      LAYER met3 ;
        RECT 1081.065000 1739.025000 1558.125000 1740.765000 ;
      LAYER met4 ;
        RECT 1081.065000 1345.985000 1082.805000 1740.765000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 2176.235000 350.985000 2177.975000 745.765000 ;
      LAYER met3 ;
        RECT 1700.915000 350.985000 2177.975000 352.725000 ;
      LAYER met3 ;
        RECT 1700.915000 744.025000 2177.975000 745.765000 ;
      LAYER met4 ;
        RECT 1700.915000 350.985000 1702.655000 745.765000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 2176.235000 848.485000 2177.975000 1243.265000 ;
      LAYER met3 ;
        RECT 1700.915000 848.485000 2177.975000 850.225000 ;
      LAYER met3 ;
        RECT 1700.915000 1241.525000 2177.975000 1243.265000 ;
      LAYER met4 ;
        RECT 1700.915000 848.485000 1702.655000 1243.265000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 2176.235000 1345.985000 2177.975000 1740.765000 ;
      LAYER met3 ;
        RECT 1700.915000 1345.985000 2177.975000 1347.725000 ;
      LAYER met3 ;
        RECT 1700.915000 1739.025000 2177.975000 1740.765000 ;
      LAYER met4 ;
        RECT 1700.915000 1345.985000 1702.655000 1740.765000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 2176.235000 1843.485000 2177.975000 2238.265000 ;
      LAYER met3 ;
        RECT 1700.915000 1843.485000 2177.975000 1845.225000 ;
      LAYER met3 ;
        RECT 1700.915000 2236.525000 2177.975000 2238.265000 ;
      LAYER met4 ;
        RECT 1700.915000 1843.485000 1702.655000 2238.265000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END vssd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 13.780000 14.060000 2212.160000 18.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780000 2875.340000 2212.160000 2879.340000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2208.160000 14.060000 2212.160000 2879.340000 ;
    END
    PORT
      LAYER met4 ;
        RECT 13.780000 14.060000 17.780000 2879.340000 ;
    END

# P/G pin shape extracted from block 'tcam_32x28'
    PORT
      LAYER met4 ;
        RECT 1581.475000 2377.035000 1583.215000 2765.015000 ;
      LAYER met4 ;
        RECT 1112.955000 2377.035000 1114.695000 2765.015000 ;
      LAYER met3 ;
        RECT 1112.955000 2377.035000 1583.215000 2378.775000 ;
      LAYER met3 ;
        RECT 1112.955000 2763.275000 1583.215000 2765.015000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2143.615000 2377.130000 2145.355000 2765.110000 ;
      LAYER met4 ;
        RECT 1675.095000 2377.130000 1676.835000 2765.110000 ;
      LAYER met3 ;
        RECT 1675.095000 2377.130000 2145.355000 2378.870000 ;
      LAYER met3 ;
        RECT 1675.095000 2763.370000 2145.355000 2765.110000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1087.285000 2338.000000 1089.285000 2800.240000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2169.225000 2338.000000 2171.225000 2800.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1087.285000 2798.240000 2171.225000 2800.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1087.285000 2338.000000 2171.225000 2340.000000 ;
    END
# end of P/G pin shape extracted from block 'tcam_32x28'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 1084.465000 740.625000 1554.725000 742.365000 ;
      LAYER met3 ;
        RECT 1084.465000 354.385000 1554.725000 356.125000 ;
      LAYER met4 ;
        RECT 1084.465000 354.385000 1086.205000 742.365000 ;
      LAYER met4 ;
        RECT 1552.985000 354.385000 1554.725000 742.365000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 1084.465000 1238.125000 1554.725000 1239.865000 ;
      LAYER met3 ;
        RECT 1084.465000 851.885000 1554.725000 853.625000 ;
      LAYER met4 ;
        RECT 1084.465000 851.885000 1086.205000 1239.865000 ;
      LAYER met4 ;
        RECT 1552.985000 851.885000 1554.725000 1239.865000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 1084.465000 2233.125000 1554.725000 2234.865000 ;
      LAYER met3 ;
        RECT 1084.465000 1846.885000 1554.725000 1848.625000 ;
      LAYER met4 ;
        RECT 1084.465000 1846.885000 1086.205000 2234.865000 ;
      LAYER met4 ;
        RECT 1552.985000 1846.885000 1554.725000 2234.865000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 1084.465000 1735.625000 1554.725000 1737.365000 ;
      LAYER met3 ;
        RECT 1084.465000 1349.385000 1554.725000 1351.125000 ;
      LAYER met4 ;
        RECT 1084.465000 1349.385000 1086.205000 1737.365000 ;
      LAYER met4 ;
        RECT 1552.985000 1349.385000 1554.725000 1737.365000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 1704.315000 740.625000 2174.575000 742.365000 ;
      LAYER met3 ;
        RECT 1704.315000 354.385000 2174.575000 356.125000 ;
      LAYER met4 ;
        RECT 1704.315000 354.385000 1706.055000 742.365000 ;
      LAYER met4 ;
        RECT 2172.835000 354.385000 2174.575000 742.365000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 1704.315000 1238.125000 2174.575000 1239.865000 ;
      LAYER met3 ;
        RECT 1704.315000 851.885000 2174.575000 853.625000 ;
      LAYER met4 ;
        RECT 1704.315000 851.885000 1706.055000 1239.865000 ;
      LAYER met4 ;
        RECT 2172.835000 851.885000 2174.575000 1239.865000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 1704.315000 1735.625000 2174.575000 1737.365000 ;
      LAYER met3 ;
        RECT 1704.315000 1349.385000 2174.575000 1351.125000 ;
      LAYER met4 ;
        RECT 1704.315000 1349.385000 1706.055000 1737.365000 ;
      LAYER met4 ;
        RECT 2172.835000 1349.385000 2174.575000 1737.365000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 1704.315000 2233.125000 2174.575000 2234.865000 ;
      LAYER met3 ;
        RECT 1704.315000 1846.885000 2174.575000 1848.625000 ;
      LAYER met4 ;
        RECT 1704.315000 1846.885000 1706.055000 2234.865000 ;
      LAYER met4 ;
        RECT 2172.835000 1846.885000 2174.575000 2234.865000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END vccd1
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 2225.940000 2895.100000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 2225.940000 2895.100000 ;
    LAYER met2 ;
      RECT 2222.610000 2894.475000 2225.940000 2895.100000 ;
      RECT 2162.510000 2894.475000 2222.190000 2895.100000 ;
      RECT 4.510000 2894.475000 63.390000 2895.100000 ;
      RECT 0.000000 2894.475000 4.090000 2895.100000 ;
      RECT 2162.510000 2894.470000 2225.940000 2894.475000 ;
      RECT 2098.910000 2894.470000 2162.090000 2895.100000 ;
      RECT 2035.310000 2894.470000 2098.490000 2895.100000 ;
      RECT 1971.710000 2894.470000 2034.890000 2895.100000 ;
      RECT 1908.110000 2894.470000 1971.290000 2895.100000 ;
      RECT 1844.510000 2894.470000 1907.690000 2895.100000 ;
      RECT 1780.910000 2894.470000 1844.090000 2895.100000 ;
      RECT 1717.310000 2894.470000 1780.490000 2895.100000 ;
      RECT 1653.710000 2894.470000 1716.890000 2895.100000 ;
      RECT 1590.110000 2894.470000 1653.290000 2895.100000 ;
      RECT 1526.510000 2894.470000 1589.690000 2895.100000 ;
      RECT 1462.910000 2894.470000 1526.090000 2895.100000 ;
      RECT 1399.310000 2894.470000 1462.490000 2895.100000 ;
      RECT 1335.710000 2894.470000 1398.890000 2895.100000 ;
      RECT 1272.110000 2894.470000 1335.290000 2895.100000 ;
      RECT 1208.510000 2894.470000 1271.690000 2895.100000 ;
      RECT 1144.910000 2894.470000 1208.090000 2895.100000 ;
      RECT 1081.310000 2894.470000 1144.490000 2895.100000 ;
      RECT 1017.710000 2894.470000 1080.890000 2895.100000 ;
      RECT 954.110000 2894.470000 1017.290000 2895.100000 ;
      RECT 890.510000 2894.470000 953.690000 2895.100000 ;
      RECT 826.910000 2894.470000 890.090000 2895.100000 ;
      RECT 763.310000 2894.470000 826.490000 2895.100000 ;
      RECT 699.710000 2894.470000 762.890000 2895.100000 ;
      RECT 636.110000 2894.470000 699.290000 2895.100000 ;
      RECT 572.510000 2894.470000 635.690000 2895.100000 ;
      RECT 508.910000 2894.470000 572.090000 2895.100000 ;
      RECT 445.310000 2894.470000 508.490000 2895.100000 ;
      RECT 381.710000 2894.470000 444.890000 2895.100000 ;
      RECT 318.110000 2894.470000 381.290000 2895.100000 ;
      RECT 254.510000 2894.470000 317.690000 2895.100000 ;
      RECT 190.910000 2894.470000 254.090000 2895.100000 ;
      RECT 127.310000 2894.470000 190.490000 2895.100000 ;
      RECT 63.810000 2894.470000 126.890000 2895.100000 ;
      RECT 0.000000 2894.470000 63.390000 2894.475000 ;
      RECT 0.000000 0.630000 2225.940000 2894.470000 ;
      RECT 2221.510000 0.625000 2225.940000 0.630000 ;
      RECT 0.000000 0.625000 4.290000 0.630000 ;
      RECT 2224.510000 0.000000 2225.940000 0.625000 ;
      RECT 2221.510000 0.000000 2224.090000 0.625000 ;
      RECT 2217.010000 0.000000 2221.090000 0.630000 ;
      RECT 2212.510000 0.000000 2216.590000 0.630000 ;
      RECT 2208.010000 0.000000 2212.090000 0.630000 ;
      RECT 2203.510000 0.000000 2207.590000 0.630000 ;
      RECT 2199.010000 0.000000 2203.090000 0.630000 ;
      RECT 2194.410000 0.000000 2198.590000 0.630000 ;
      RECT 2189.910000 0.000000 2193.990000 0.630000 ;
      RECT 2185.410000 0.000000 2189.490000 0.630000 ;
      RECT 2180.910000 0.000000 2184.990000 0.630000 ;
      RECT 2176.410000 0.000000 2180.490000 0.630000 ;
      RECT 2171.910000 0.000000 2175.990000 0.630000 ;
      RECT 2167.410000 0.000000 2171.490000 0.630000 ;
      RECT 2162.810000 0.000000 2166.990000 0.630000 ;
      RECT 2158.310000 0.000000 2162.390000 0.630000 ;
      RECT 2153.810000 0.000000 2157.890000 0.630000 ;
      RECT 2149.310000 0.000000 2153.390000 0.630000 ;
      RECT 2144.810000 0.000000 2148.890000 0.630000 ;
      RECT 2140.310000 0.000000 2144.390000 0.630000 ;
      RECT 2135.710000 0.000000 2139.890000 0.630000 ;
      RECT 2131.210000 0.000000 2135.290000 0.630000 ;
      RECT 2126.710000 0.000000 2130.790000 0.630000 ;
      RECT 2122.210000 0.000000 2126.290000 0.630000 ;
      RECT 2117.710000 0.000000 2121.790000 0.630000 ;
      RECT 2113.210000 0.000000 2117.290000 0.630000 ;
      RECT 2108.710000 0.000000 2112.790000 0.630000 ;
      RECT 2104.110000 0.000000 2108.290000 0.630000 ;
      RECT 2099.610000 0.000000 2103.690000 0.630000 ;
      RECT 2095.110000 0.000000 2099.190000 0.630000 ;
      RECT 2090.610000 0.000000 2094.690000 0.630000 ;
      RECT 2086.110000 0.000000 2090.190000 0.630000 ;
      RECT 2081.610000 0.000000 2085.690000 0.630000 ;
      RECT 2077.110000 0.000000 2081.190000 0.630000 ;
      RECT 2072.510000 0.000000 2076.690000 0.630000 ;
      RECT 2068.010000 0.000000 2072.090000 0.630000 ;
      RECT 2063.510000 0.000000 2067.590000 0.630000 ;
      RECT 2059.010000 0.000000 2063.090000 0.630000 ;
      RECT 2054.510000 0.000000 2058.590000 0.630000 ;
      RECT 2050.010000 0.000000 2054.090000 0.630000 ;
      RECT 2045.410000 0.000000 2049.590000 0.630000 ;
      RECT 2040.910000 0.000000 2044.990000 0.630000 ;
      RECT 2036.410000 0.000000 2040.490000 0.630000 ;
      RECT 2031.910000 0.000000 2035.990000 0.630000 ;
      RECT 2027.410000 0.000000 2031.490000 0.630000 ;
      RECT 2022.910000 0.000000 2026.990000 0.630000 ;
      RECT 2018.410000 0.000000 2022.490000 0.630000 ;
      RECT 2013.810000 0.000000 2017.990000 0.630000 ;
      RECT 2009.310000 0.000000 2013.390000 0.630000 ;
      RECT 2004.810000 0.000000 2008.890000 0.630000 ;
      RECT 2000.310000 0.000000 2004.390000 0.630000 ;
      RECT 1995.810000 0.000000 1999.890000 0.630000 ;
      RECT 1991.310000 0.000000 1995.390000 0.630000 ;
      RECT 1986.810000 0.000000 1990.890000 0.630000 ;
      RECT 1982.210000 0.000000 1986.390000 0.630000 ;
      RECT 1977.710000 0.000000 1981.790000 0.630000 ;
      RECT 1973.210000 0.000000 1977.290000 0.630000 ;
      RECT 1968.710000 0.000000 1972.790000 0.630000 ;
      RECT 1964.210000 0.000000 1968.290000 0.630000 ;
      RECT 1959.710000 0.000000 1963.790000 0.630000 ;
      RECT 1955.110000 0.000000 1959.290000 0.630000 ;
      RECT 1950.610000 0.000000 1954.690000 0.630000 ;
      RECT 1946.110000 0.000000 1950.190000 0.630000 ;
      RECT 1941.610000 0.000000 1945.690000 0.630000 ;
      RECT 1937.110000 0.000000 1941.190000 0.630000 ;
      RECT 1932.610000 0.000000 1936.690000 0.630000 ;
      RECT 1928.110000 0.000000 1932.190000 0.630000 ;
      RECT 1923.510000 0.000000 1927.690000 0.630000 ;
      RECT 1919.010000 0.000000 1923.090000 0.630000 ;
      RECT 1914.510000 0.000000 1918.590000 0.630000 ;
      RECT 1910.010000 0.000000 1914.090000 0.630000 ;
      RECT 1905.510000 0.000000 1909.590000 0.630000 ;
      RECT 1901.010000 0.000000 1905.090000 0.630000 ;
      RECT 1896.510000 0.000000 1900.590000 0.630000 ;
      RECT 1891.910000 0.000000 1896.090000 0.630000 ;
      RECT 1887.410000 0.000000 1891.490000 0.630000 ;
      RECT 1882.910000 0.000000 1886.990000 0.630000 ;
      RECT 1878.410000 0.000000 1882.490000 0.630000 ;
      RECT 1873.910000 0.000000 1877.990000 0.630000 ;
      RECT 1869.410000 0.000000 1873.490000 0.630000 ;
      RECT 1864.810000 0.000000 1868.990000 0.630000 ;
      RECT 1860.310000 0.000000 1864.390000 0.630000 ;
      RECT 1855.810000 0.000000 1859.890000 0.630000 ;
      RECT 1851.310000 0.000000 1855.390000 0.630000 ;
      RECT 1846.810000 0.000000 1850.890000 0.630000 ;
      RECT 1842.310000 0.000000 1846.390000 0.630000 ;
      RECT 1837.810000 0.000000 1841.890000 0.630000 ;
      RECT 1833.210000 0.000000 1837.390000 0.630000 ;
      RECT 1828.710000 0.000000 1832.790000 0.630000 ;
      RECT 1824.210000 0.000000 1828.290000 0.630000 ;
      RECT 1819.710000 0.000000 1823.790000 0.630000 ;
      RECT 1815.210000 0.000000 1819.290000 0.630000 ;
      RECT 1810.710000 0.000000 1814.790000 0.630000 ;
      RECT 1806.210000 0.000000 1810.290000 0.630000 ;
      RECT 1801.610000 0.000000 1805.790000 0.630000 ;
      RECT 1797.110000 0.000000 1801.190000 0.630000 ;
      RECT 1792.610000 0.000000 1796.690000 0.630000 ;
      RECT 1788.110000 0.000000 1792.190000 0.630000 ;
      RECT 1783.610000 0.000000 1787.690000 0.630000 ;
      RECT 1779.110000 0.000000 1783.190000 0.630000 ;
      RECT 1774.510000 0.000000 1778.690000 0.630000 ;
      RECT 1770.010000 0.000000 1774.090000 0.630000 ;
      RECT 1765.510000 0.000000 1769.590000 0.630000 ;
      RECT 1761.010000 0.000000 1765.090000 0.630000 ;
      RECT 1756.510000 0.000000 1760.590000 0.630000 ;
      RECT 1752.010000 0.000000 1756.090000 0.630000 ;
      RECT 1747.510000 0.000000 1751.590000 0.630000 ;
      RECT 1742.910000 0.000000 1747.090000 0.630000 ;
      RECT 1738.410000 0.000000 1742.490000 0.630000 ;
      RECT 1733.910000 0.000000 1737.990000 0.630000 ;
      RECT 1729.410000 0.000000 1733.490000 0.630000 ;
      RECT 1724.910000 0.000000 1728.990000 0.630000 ;
      RECT 1720.410000 0.000000 1724.490000 0.630000 ;
      RECT 1715.910000 0.000000 1719.990000 0.630000 ;
      RECT 1711.310000 0.000000 1715.490000 0.630000 ;
      RECT 1706.810000 0.000000 1710.890000 0.630000 ;
      RECT 1702.310000 0.000000 1706.390000 0.630000 ;
      RECT 1697.810000 0.000000 1701.890000 0.630000 ;
      RECT 1693.310000 0.000000 1697.390000 0.630000 ;
      RECT 1688.810000 0.000000 1692.890000 0.630000 ;
      RECT 1684.210000 0.000000 1688.390000 0.630000 ;
      RECT 1679.710000 0.000000 1683.790000 0.630000 ;
      RECT 1675.210000 0.000000 1679.290000 0.630000 ;
      RECT 1670.710000 0.000000 1674.790000 0.630000 ;
      RECT 1666.210000 0.000000 1670.290000 0.630000 ;
      RECT 1661.710000 0.000000 1665.790000 0.630000 ;
      RECT 1657.210000 0.000000 1661.290000 0.630000 ;
      RECT 1652.610000 0.000000 1656.790000 0.630000 ;
      RECT 1648.110000 0.000000 1652.190000 0.630000 ;
      RECT 1643.610000 0.000000 1647.690000 0.630000 ;
      RECT 1639.110000 0.000000 1643.190000 0.630000 ;
      RECT 1634.610000 0.000000 1638.690000 0.630000 ;
      RECT 1630.110000 0.000000 1634.190000 0.630000 ;
      RECT 1625.610000 0.000000 1629.690000 0.630000 ;
      RECT 1621.010000 0.000000 1625.190000 0.630000 ;
      RECT 1616.510000 0.000000 1620.590000 0.630000 ;
      RECT 1612.010000 0.000000 1616.090000 0.630000 ;
      RECT 1607.510000 0.000000 1611.590000 0.630000 ;
      RECT 1603.010000 0.000000 1607.090000 0.630000 ;
      RECT 1598.510000 0.000000 1602.590000 0.630000 ;
      RECT 1593.910000 0.000000 1598.090000 0.630000 ;
      RECT 1589.410000 0.000000 1593.490000 0.630000 ;
      RECT 1584.910000 0.000000 1588.990000 0.630000 ;
      RECT 1580.410000 0.000000 1584.490000 0.630000 ;
      RECT 1575.910000 0.000000 1579.990000 0.630000 ;
      RECT 1571.410000 0.000000 1575.490000 0.630000 ;
      RECT 1566.910000 0.000000 1570.990000 0.630000 ;
      RECT 1562.310000 0.000000 1566.490000 0.630000 ;
      RECT 1557.810000 0.000000 1561.890000 0.630000 ;
      RECT 1553.310000 0.000000 1557.390000 0.630000 ;
      RECT 1548.810000 0.000000 1552.890000 0.630000 ;
      RECT 1544.310000 0.000000 1548.390000 0.630000 ;
      RECT 1539.810000 0.000000 1543.890000 0.630000 ;
      RECT 1535.310000 0.000000 1539.390000 0.630000 ;
      RECT 1530.710000 0.000000 1534.890000 0.630000 ;
      RECT 1526.210000 0.000000 1530.290000 0.630000 ;
      RECT 1521.710000 0.000000 1525.790000 0.630000 ;
      RECT 1517.210000 0.000000 1521.290000 0.630000 ;
      RECT 1512.710000 0.000000 1516.790000 0.630000 ;
      RECT 1508.210000 0.000000 1512.290000 0.630000 ;
      RECT 1503.610000 0.000000 1507.790000 0.630000 ;
      RECT 1499.110000 0.000000 1503.190000 0.630000 ;
      RECT 1494.610000 0.000000 1498.690000 0.630000 ;
      RECT 1490.110000 0.000000 1494.190000 0.630000 ;
      RECT 1485.610000 0.000000 1489.690000 0.630000 ;
      RECT 1481.110000 0.000000 1485.190000 0.630000 ;
      RECT 1476.610000 0.000000 1480.690000 0.630000 ;
      RECT 1472.010000 0.000000 1476.190000 0.630000 ;
      RECT 1467.510000 0.000000 1471.590000 0.630000 ;
      RECT 1463.010000 0.000000 1467.090000 0.630000 ;
      RECT 1458.510000 0.000000 1462.590000 0.630000 ;
      RECT 1454.010000 0.000000 1458.090000 0.630000 ;
      RECT 1449.510000 0.000000 1453.590000 0.630000 ;
      RECT 1445.010000 0.000000 1449.090000 0.630000 ;
      RECT 1440.410000 0.000000 1444.590000 0.630000 ;
      RECT 1435.910000 0.000000 1439.990000 0.630000 ;
      RECT 1431.410000 0.000000 1435.490000 0.630000 ;
      RECT 1426.910000 0.000000 1430.990000 0.630000 ;
      RECT 1422.410000 0.000000 1426.490000 0.630000 ;
      RECT 1417.910000 0.000000 1421.990000 0.630000 ;
      RECT 1413.310000 0.000000 1417.490000 0.630000 ;
      RECT 1408.810000 0.000000 1412.890000 0.630000 ;
      RECT 1404.310000 0.000000 1408.390000 0.630000 ;
      RECT 1399.810000 0.000000 1403.890000 0.630000 ;
      RECT 1395.310000 0.000000 1399.390000 0.630000 ;
      RECT 1390.810000 0.000000 1394.890000 0.630000 ;
      RECT 1386.310000 0.000000 1390.390000 0.630000 ;
      RECT 1381.710000 0.000000 1385.890000 0.630000 ;
      RECT 1377.210000 0.000000 1381.290000 0.630000 ;
      RECT 1372.710000 0.000000 1376.790000 0.630000 ;
      RECT 1368.210000 0.000000 1372.290000 0.630000 ;
      RECT 1363.710000 0.000000 1367.790000 0.630000 ;
      RECT 1359.210000 0.000000 1363.290000 0.630000 ;
      RECT 1354.710000 0.000000 1358.790000 0.630000 ;
      RECT 1350.110000 0.000000 1354.290000 0.630000 ;
      RECT 1345.610000 0.000000 1349.690000 0.630000 ;
      RECT 1341.110000 0.000000 1345.190000 0.630000 ;
      RECT 1336.610000 0.000000 1340.690000 0.630000 ;
      RECT 1332.110000 0.000000 1336.190000 0.630000 ;
      RECT 1327.610000 0.000000 1331.690000 0.630000 ;
      RECT 1323.010000 0.000000 1327.190000 0.630000 ;
      RECT 1318.510000 0.000000 1322.590000 0.630000 ;
      RECT 1314.010000 0.000000 1318.090000 0.630000 ;
      RECT 1309.510000 0.000000 1313.590000 0.630000 ;
      RECT 1305.010000 0.000000 1309.090000 0.630000 ;
      RECT 1300.510000 0.000000 1304.590000 0.630000 ;
      RECT 1296.010000 0.000000 1300.090000 0.630000 ;
      RECT 1291.410000 0.000000 1295.590000 0.630000 ;
      RECT 1286.910000 0.000000 1290.990000 0.630000 ;
      RECT 1282.410000 0.000000 1286.490000 0.630000 ;
      RECT 1277.910000 0.000000 1281.990000 0.630000 ;
      RECT 1273.410000 0.000000 1277.490000 0.630000 ;
      RECT 1268.910000 0.000000 1272.990000 0.630000 ;
      RECT 1264.410000 0.000000 1268.490000 0.630000 ;
      RECT 1259.810000 0.000000 1263.990000 0.630000 ;
      RECT 1255.310000 0.000000 1259.390000 0.630000 ;
      RECT 1250.810000 0.000000 1254.890000 0.630000 ;
      RECT 1246.310000 0.000000 1250.390000 0.630000 ;
      RECT 1241.810000 0.000000 1245.890000 0.630000 ;
      RECT 1237.310000 0.000000 1241.390000 0.630000 ;
      RECT 1232.710000 0.000000 1236.890000 0.630000 ;
      RECT 1228.210000 0.000000 1232.290000 0.630000 ;
      RECT 1223.710000 0.000000 1227.790000 0.630000 ;
      RECT 1219.210000 0.000000 1223.290000 0.630000 ;
      RECT 1214.710000 0.000000 1218.790000 0.630000 ;
      RECT 1210.210000 0.000000 1214.290000 0.630000 ;
      RECT 1205.710000 0.000000 1209.790000 0.630000 ;
      RECT 1201.110000 0.000000 1205.290000 0.630000 ;
      RECT 1196.610000 0.000000 1200.690000 0.630000 ;
      RECT 1192.110000 0.000000 1196.190000 0.630000 ;
      RECT 1187.610000 0.000000 1191.690000 0.630000 ;
      RECT 1183.110000 0.000000 1187.190000 0.630000 ;
      RECT 1178.610000 0.000000 1182.690000 0.630000 ;
      RECT 1174.110000 0.000000 1178.190000 0.630000 ;
      RECT 1169.510000 0.000000 1173.690000 0.630000 ;
      RECT 1165.010000 0.000000 1169.090000 0.630000 ;
      RECT 1160.510000 0.000000 1164.590000 0.630000 ;
      RECT 1156.010000 0.000000 1160.090000 0.630000 ;
      RECT 1151.510000 0.000000 1155.590000 0.630000 ;
      RECT 1147.010000 0.000000 1151.090000 0.630000 ;
      RECT 1142.410000 0.000000 1146.590000 0.630000 ;
      RECT 1137.910000 0.000000 1141.990000 0.630000 ;
      RECT 1133.410000 0.000000 1137.490000 0.630000 ;
      RECT 1128.910000 0.000000 1132.990000 0.630000 ;
      RECT 1124.410000 0.000000 1128.490000 0.630000 ;
      RECT 1119.910000 0.000000 1123.990000 0.630000 ;
      RECT 1115.410000 0.000000 1119.490000 0.630000 ;
      RECT 1110.810000 0.000000 1114.990000 0.630000 ;
      RECT 1106.310000 0.000000 1110.390000 0.630000 ;
      RECT 1101.810000 0.000000 1105.890000 0.630000 ;
      RECT 1097.310000 0.000000 1101.390000 0.630000 ;
      RECT 1092.810000 0.000000 1096.890000 0.630000 ;
      RECT 1088.310000 0.000000 1092.390000 0.630000 ;
      RECT 1083.810000 0.000000 1087.890000 0.630000 ;
      RECT 1079.210000 0.000000 1083.390000 0.630000 ;
      RECT 1074.710000 0.000000 1078.790000 0.630000 ;
      RECT 1070.210000 0.000000 1074.290000 0.630000 ;
      RECT 1065.710000 0.000000 1069.790000 0.630000 ;
      RECT 1061.210000 0.000000 1065.290000 0.630000 ;
      RECT 1056.710000 0.000000 1060.790000 0.630000 ;
      RECT 1052.110000 0.000000 1056.290000 0.630000 ;
      RECT 1047.610000 0.000000 1051.690000 0.630000 ;
      RECT 1043.110000 0.000000 1047.190000 0.630000 ;
      RECT 1038.610000 0.000000 1042.690000 0.630000 ;
      RECT 1034.110000 0.000000 1038.190000 0.630000 ;
      RECT 1029.610000 0.000000 1033.690000 0.630000 ;
      RECT 1025.110000 0.000000 1029.190000 0.630000 ;
      RECT 1020.510000 0.000000 1024.690000 0.630000 ;
      RECT 1016.010000 0.000000 1020.090000 0.630000 ;
      RECT 1011.510000 0.000000 1015.590000 0.630000 ;
      RECT 1007.010000 0.000000 1011.090000 0.630000 ;
      RECT 1002.510000 0.000000 1006.590000 0.630000 ;
      RECT 998.010000 0.000000 1002.090000 0.630000 ;
      RECT 993.510000 0.000000 997.590000 0.630000 ;
      RECT 988.910000 0.000000 993.090000 0.630000 ;
      RECT 984.410000 0.000000 988.490000 0.630000 ;
      RECT 979.910000 0.000000 983.990000 0.630000 ;
      RECT 975.410000 0.000000 979.490000 0.630000 ;
      RECT 970.910000 0.000000 974.990000 0.630000 ;
      RECT 966.410000 0.000000 970.490000 0.630000 ;
      RECT 961.810000 0.000000 965.990000 0.630000 ;
      RECT 957.310000 0.000000 961.390000 0.630000 ;
      RECT 952.810000 0.000000 956.890000 0.630000 ;
      RECT 948.310000 0.000000 952.390000 0.630000 ;
      RECT 943.810000 0.000000 947.890000 0.630000 ;
      RECT 939.310000 0.000000 943.390000 0.630000 ;
      RECT 934.810000 0.000000 938.890000 0.630000 ;
      RECT 930.210000 0.000000 934.390000 0.630000 ;
      RECT 925.710000 0.000000 929.790000 0.630000 ;
      RECT 921.210000 0.000000 925.290000 0.630000 ;
      RECT 916.710000 0.000000 920.790000 0.630000 ;
      RECT 912.210000 0.000000 916.290000 0.630000 ;
      RECT 907.710000 0.000000 911.790000 0.630000 ;
      RECT 903.210000 0.000000 907.290000 0.630000 ;
      RECT 898.610000 0.000000 902.790000 0.630000 ;
      RECT 894.110000 0.000000 898.190000 0.630000 ;
      RECT 889.610000 0.000000 893.690000 0.630000 ;
      RECT 885.110000 0.000000 889.190000 0.630000 ;
      RECT 880.610000 0.000000 884.690000 0.630000 ;
      RECT 876.110000 0.000000 880.190000 0.630000 ;
      RECT 871.510000 0.000000 875.690000 0.630000 ;
      RECT 867.010000 0.000000 871.090000 0.630000 ;
      RECT 862.510000 0.000000 866.590000 0.630000 ;
      RECT 858.010000 0.000000 862.090000 0.630000 ;
      RECT 853.510000 0.000000 857.590000 0.630000 ;
      RECT 849.010000 0.000000 853.090000 0.630000 ;
      RECT 844.510000 0.000000 848.590000 0.630000 ;
      RECT 839.910000 0.000000 844.090000 0.630000 ;
      RECT 835.410000 0.000000 839.490000 0.630000 ;
      RECT 830.910000 0.000000 834.990000 0.630000 ;
      RECT 826.410000 0.000000 830.490000 0.630000 ;
      RECT 821.910000 0.000000 825.990000 0.630000 ;
      RECT 817.410000 0.000000 821.490000 0.630000 ;
      RECT 812.910000 0.000000 816.990000 0.630000 ;
      RECT 808.310000 0.000000 812.490000 0.630000 ;
      RECT 803.810000 0.000000 807.890000 0.630000 ;
      RECT 799.310000 0.000000 803.390000 0.630000 ;
      RECT 794.810000 0.000000 798.890000 0.630000 ;
      RECT 790.310000 0.000000 794.390000 0.630000 ;
      RECT 785.810000 0.000000 789.890000 0.630000 ;
      RECT 781.210000 0.000000 785.390000 0.630000 ;
      RECT 776.710000 0.000000 780.790000 0.630000 ;
      RECT 772.210000 0.000000 776.290000 0.630000 ;
      RECT 767.710000 0.000000 771.790000 0.630000 ;
      RECT 763.210000 0.000000 767.290000 0.630000 ;
      RECT 758.710000 0.000000 762.790000 0.630000 ;
      RECT 754.210000 0.000000 758.290000 0.630000 ;
      RECT 749.610000 0.000000 753.790000 0.630000 ;
      RECT 745.110000 0.000000 749.190000 0.630000 ;
      RECT 740.610000 0.000000 744.690000 0.630000 ;
      RECT 736.110000 0.000000 740.190000 0.630000 ;
      RECT 731.610000 0.000000 735.690000 0.630000 ;
      RECT 727.110000 0.000000 731.190000 0.630000 ;
      RECT 722.610000 0.000000 726.690000 0.630000 ;
      RECT 718.010000 0.000000 722.190000 0.630000 ;
      RECT 713.510000 0.000000 717.590000 0.630000 ;
      RECT 709.010000 0.000000 713.090000 0.630000 ;
      RECT 704.510000 0.000000 708.590000 0.630000 ;
      RECT 700.010000 0.000000 704.090000 0.630000 ;
      RECT 695.510000 0.000000 699.590000 0.630000 ;
      RECT 690.910000 0.000000 695.090000 0.630000 ;
      RECT 686.410000 0.000000 690.490000 0.630000 ;
      RECT 681.910000 0.000000 685.990000 0.630000 ;
      RECT 677.410000 0.000000 681.490000 0.630000 ;
      RECT 672.910000 0.000000 676.990000 0.630000 ;
      RECT 668.410000 0.000000 672.490000 0.630000 ;
      RECT 663.910000 0.000000 667.990000 0.630000 ;
      RECT 659.310000 0.000000 663.490000 0.630000 ;
      RECT 654.810000 0.000000 658.890000 0.630000 ;
      RECT 650.310000 0.000000 654.390000 0.630000 ;
      RECT 645.810000 0.000000 649.890000 0.630000 ;
      RECT 641.310000 0.000000 645.390000 0.630000 ;
      RECT 636.810000 0.000000 640.890000 0.630000 ;
      RECT 632.310000 0.000000 636.390000 0.630000 ;
      RECT 627.710000 0.000000 631.890000 0.630000 ;
      RECT 623.210000 0.000000 627.290000 0.630000 ;
      RECT 618.710000 0.000000 622.790000 0.630000 ;
      RECT 614.210000 0.000000 618.290000 0.630000 ;
      RECT 609.710000 0.000000 613.790000 0.630000 ;
      RECT 605.210000 0.000000 609.290000 0.630000 ;
      RECT 600.610000 0.000000 604.790000 0.630000 ;
      RECT 596.110000 0.000000 600.190000 0.630000 ;
      RECT 591.610000 0.000000 595.690000 0.630000 ;
      RECT 587.110000 0.000000 591.190000 0.630000 ;
      RECT 582.610000 0.000000 586.690000 0.630000 ;
      RECT 578.110000 0.000000 582.190000 0.630000 ;
      RECT 573.610000 0.000000 577.690000 0.630000 ;
      RECT 569.010000 0.000000 573.190000 0.630000 ;
      RECT 564.510000 0.000000 568.590000 0.630000 ;
      RECT 560.010000 0.000000 564.090000 0.630000 ;
      RECT 555.510000 0.000000 559.590000 0.630000 ;
      RECT 551.010000 0.000000 555.090000 0.630000 ;
      RECT 546.510000 0.000000 550.590000 0.630000 ;
      RECT 542.010000 0.000000 546.090000 0.630000 ;
      RECT 537.410000 0.000000 541.590000 0.630000 ;
      RECT 532.910000 0.000000 536.990000 0.630000 ;
      RECT 528.410000 0.000000 532.490000 0.630000 ;
      RECT 523.910000 0.000000 527.990000 0.630000 ;
      RECT 519.410000 0.000000 523.490000 0.630000 ;
      RECT 514.910000 0.000000 518.990000 0.630000 ;
      RECT 510.310000 0.000000 514.490000 0.630000 ;
      RECT 505.810000 0.000000 509.890000 0.630000 ;
      RECT 501.310000 0.000000 505.390000 0.630000 ;
      RECT 496.810000 0.000000 500.890000 0.630000 ;
      RECT 492.310000 0.000000 496.390000 0.630000 ;
      RECT 487.810000 0.000000 491.890000 0.630000 ;
      RECT 483.310000 0.000000 487.390000 0.630000 ;
      RECT 478.710000 0.000000 482.890000 0.630000 ;
      RECT 474.210000 0.000000 478.290000 0.630000 ;
      RECT 469.710000 0.000000 473.790000 0.630000 ;
      RECT 465.210000 0.000000 469.290000 0.630000 ;
      RECT 460.710000 0.000000 464.790000 0.630000 ;
      RECT 456.210000 0.000000 460.290000 0.630000 ;
      RECT 451.710000 0.000000 455.790000 0.630000 ;
      RECT 447.110000 0.000000 451.290000 0.630000 ;
      RECT 442.610000 0.000000 446.690000 0.630000 ;
      RECT 438.110000 0.000000 442.190000 0.630000 ;
      RECT 433.610000 0.000000 437.690000 0.630000 ;
      RECT 429.110000 0.000000 433.190000 0.630000 ;
      RECT 424.610000 0.000000 428.690000 0.630000 ;
      RECT 420.010000 0.000000 424.190000 0.630000 ;
      RECT 415.510000 0.000000 419.590000 0.630000 ;
      RECT 411.010000 0.000000 415.090000 0.630000 ;
      RECT 406.510000 0.000000 410.590000 0.630000 ;
      RECT 402.010000 0.000000 406.090000 0.630000 ;
      RECT 397.510000 0.000000 401.590000 0.630000 ;
      RECT 393.010000 0.000000 397.090000 0.630000 ;
      RECT 388.410000 0.000000 392.590000 0.630000 ;
      RECT 383.910000 0.000000 387.990000 0.630000 ;
      RECT 379.410000 0.000000 383.490000 0.630000 ;
      RECT 374.910000 0.000000 378.990000 0.630000 ;
      RECT 370.410000 0.000000 374.490000 0.630000 ;
      RECT 365.910000 0.000000 369.990000 0.630000 ;
      RECT 361.410000 0.000000 365.490000 0.630000 ;
      RECT 356.810000 0.000000 360.990000 0.630000 ;
      RECT 352.310000 0.000000 356.390000 0.630000 ;
      RECT 347.810000 0.000000 351.890000 0.630000 ;
      RECT 343.310000 0.000000 347.390000 0.630000 ;
      RECT 338.810000 0.000000 342.890000 0.630000 ;
      RECT 334.310000 0.000000 338.390000 0.630000 ;
      RECT 329.710000 0.000000 333.890000 0.630000 ;
      RECT 325.210000 0.000000 329.290000 0.630000 ;
      RECT 320.710000 0.000000 324.790000 0.630000 ;
      RECT 316.210000 0.000000 320.290000 0.630000 ;
      RECT 311.710000 0.000000 315.790000 0.630000 ;
      RECT 307.210000 0.000000 311.290000 0.630000 ;
      RECT 302.710000 0.000000 306.790000 0.630000 ;
      RECT 298.110000 0.000000 302.290000 0.630000 ;
      RECT 293.610000 0.000000 297.690000 0.630000 ;
      RECT 289.110000 0.000000 293.190000 0.630000 ;
      RECT 284.610000 0.000000 288.690000 0.630000 ;
      RECT 280.110000 0.000000 284.190000 0.630000 ;
      RECT 275.610000 0.000000 279.690000 0.630000 ;
      RECT 271.110000 0.000000 275.190000 0.630000 ;
      RECT 266.510000 0.000000 270.690000 0.630000 ;
      RECT 262.010000 0.000000 266.090000 0.630000 ;
      RECT 257.510000 0.000000 261.590000 0.630000 ;
      RECT 253.010000 0.000000 257.090000 0.630000 ;
      RECT 248.510000 0.000000 252.590000 0.630000 ;
      RECT 244.010000 0.000000 248.090000 0.630000 ;
      RECT 239.410000 0.000000 243.590000 0.630000 ;
      RECT 234.910000 0.000000 238.990000 0.630000 ;
      RECT 230.410000 0.000000 234.490000 0.630000 ;
      RECT 225.910000 0.000000 229.990000 0.630000 ;
      RECT 221.410000 0.000000 225.490000 0.630000 ;
      RECT 216.910000 0.000000 220.990000 0.630000 ;
      RECT 212.410000 0.000000 216.490000 0.630000 ;
      RECT 207.810000 0.000000 211.990000 0.630000 ;
      RECT 203.310000 0.000000 207.390000 0.630000 ;
      RECT 198.810000 0.000000 202.890000 0.630000 ;
      RECT 194.310000 0.000000 198.390000 0.630000 ;
      RECT 189.810000 0.000000 193.890000 0.630000 ;
      RECT 185.310000 0.000000 189.390000 0.630000 ;
      RECT 180.810000 0.000000 184.890000 0.630000 ;
      RECT 176.210000 0.000000 180.390000 0.630000 ;
      RECT 171.710000 0.000000 175.790000 0.630000 ;
      RECT 167.210000 0.000000 171.290000 0.630000 ;
      RECT 162.710000 0.000000 166.790000 0.630000 ;
      RECT 158.210000 0.000000 162.290000 0.630000 ;
      RECT 153.710000 0.000000 157.790000 0.630000 ;
      RECT 149.110000 0.000000 153.290000 0.630000 ;
      RECT 144.610000 0.000000 148.690000 0.630000 ;
      RECT 140.110000 0.000000 144.190000 0.630000 ;
      RECT 135.610000 0.000000 139.690000 0.630000 ;
      RECT 131.110000 0.000000 135.190000 0.630000 ;
      RECT 126.610000 0.000000 130.690000 0.630000 ;
      RECT 122.110000 0.000000 126.190000 0.630000 ;
      RECT 117.510000 0.000000 121.690000 0.630000 ;
      RECT 113.010000 0.000000 117.090000 0.630000 ;
      RECT 108.510000 0.000000 112.590000 0.630000 ;
      RECT 104.010000 0.000000 108.090000 0.630000 ;
      RECT 99.510000 0.000000 103.590000 0.630000 ;
      RECT 95.010000 0.000000 99.090000 0.630000 ;
      RECT 90.510000 0.000000 94.590000 0.630000 ;
      RECT 85.910000 0.000000 90.090000 0.630000 ;
      RECT 81.410000 0.000000 85.490000 0.630000 ;
      RECT 76.910000 0.000000 80.990000 0.630000 ;
      RECT 72.410000 0.000000 76.490000 0.630000 ;
      RECT 67.910000 0.000000 71.990000 0.630000 ;
      RECT 63.410000 0.000000 67.490000 0.630000 ;
      RECT 58.810000 0.000000 62.990000 0.630000 ;
      RECT 54.310000 0.000000 58.390000 0.630000 ;
      RECT 49.810000 0.000000 53.890000 0.630000 ;
      RECT 45.310000 0.000000 49.390000 0.630000 ;
      RECT 40.810000 0.000000 44.890000 0.630000 ;
      RECT 36.310000 0.000000 40.390000 0.630000 ;
      RECT 31.810000 0.000000 35.890000 0.630000 ;
      RECT 27.210000 0.000000 31.390000 0.630000 ;
      RECT 22.710000 0.000000 26.790000 0.630000 ;
      RECT 18.210000 0.000000 22.290000 0.630000 ;
      RECT 13.710000 0.000000 17.790000 0.630000 ;
      RECT 9.210000 0.000000 13.290000 0.630000 ;
      RECT 4.710000 0.000000 8.790000 0.630000 ;
      RECT 2.710000 0.000000 4.290000 0.625000 ;
      RECT 0.000000 0.000000 2.290000 0.625000 ;
    LAYER met3 ;
      RECT 0.000000 2885.540000 2225.940000 2895.100000 ;
      RECT 2218.360000 2884.295000 2225.940000 2885.540000 ;
      RECT 0.000000 2883.710000 7.580000 2885.540000 ;
      RECT 2218.360000 2883.395000 2224.840000 2884.295000 ;
      RECT 1.100000 2882.810000 7.580000 2883.710000 ;
      RECT 2218.360000 2880.740000 2225.940000 2883.395000 ;
      RECT 0.000000 2880.740000 7.580000 2882.810000 ;
      RECT 0.000000 2879.740000 2225.940000 2880.740000 ;
      RECT 2212.560000 2874.940000 2225.940000 2879.740000 ;
      RECT 0.000000 2874.940000 13.380000 2879.740000 ;
      RECT 0.000000 2832.060000 2225.940000 2874.940000 ;
      RECT 1.100000 2831.160000 2225.940000 2832.060000 ;
      RECT 0.000000 2831.080000 2225.940000 2831.160000 ;
      RECT 0.000000 2830.180000 2224.840000 2831.080000 ;
      RECT 0.000000 2777.670000 2225.940000 2830.180000 ;
      RECT 1.100000 2776.770000 2225.940000 2777.670000 ;
      RECT 0.000000 2775.615000 2225.940000 2776.770000 ;
      RECT 0.000000 2774.715000 2224.840000 2775.615000 ;
      RECT 0.000000 2723.185000 2225.940000 2774.715000 ;
      RECT 1.100000 2722.285000 2225.940000 2723.185000 ;
      RECT 0.000000 2720.050000 2225.940000 2722.285000 ;
      RECT 0.000000 2719.150000 2224.840000 2720.050000 ;
      RECT 0.000000 2668.695000 2225.940000 2719.150000 ;
      RECT 1.100000 2667.795000 2225.940000 2668.695000 ;
      RECT 0.000000 2664.580000 2225.940000 2667.795000 ;
      RECT 0.000000 2663.680000 2224.840000 2664.580000 ;
      RECT 0.000000 2614.305000 2225.940000 2663.680000 ;
      RECT 1.100000 2613.405000 2225.940000 2614.305000 ;
      RECT 0.000000 2609.015000 2225.940000 2613.405000 ;
      RECT 0.000000 2608.115000 2224.840000 2609.015000 ;
      RECT 0.000000 2559.820000 2225.940000 2608.115000 ;
      RECT 1.100000 2558.920000 2225.940000 2559.820000 ;
      RECT 0.000000 2553.545000 2225.940000 2558.920000 ;
      RECT 0.000000 2552.645000 2224.840000 2553.545000 ;
      RECT 0.000000 2505.330000 2225.940000 2552.645000 ;
      RECT 1.100000 2504.430000 2225.940000 2505.330000 ;
      RECT 0.000000 2498.080000 2225.940000 2504.430000 ;
      RECT 0.000000 2497.180000 2224.840000 2498.080000 ;
      RECT 0.000000 2450.940000 2225.940000 2497.180000 ;
      RECT 1.100000 2450.040000 2225.940000 2450.940000 ;
      RECT 0.000000 2442.510000 2225.940000 2450.040000 ;
      RECT 0.000000 2441.610000 2224.840000 2442.510000 ;
      RECT 0.000000 2396.450000 2225.940000 2441.610000 ;
      RECT 1.100000 2395.550000 2225.940000 2396.450000 ;
      RECT 0.000000 2387.045000 2225.940000 2395.550000 ;
      RECT 0.000000 2386.145000 2224.840000 2387.045000 ;
      RECT 0.000000 2341.965000 2225.940000 2386.145000 ;
      RECT 1.100000 2341.065000 2225.940000 2341.965000 ;
      RECT 0.000000 2331.575000 2225.940000 2341.065000 ;
      RECT 0.000000 2330.675000 2224.840000 2331.575000 ;
      RECT 0.000000 2287.575000 2225.940000 2330.675000 ;
      RECT 1.100000 2286.675000 2225.940000 2287.575000 ;
      RECT 0.000000 2276.010000 2225.940000 2286.675000 ;
      RECT 0.000000 2275.110000 2224.840000 2276.010000 ;
      RECT 0.000000 2233.085000 2225.940000 2275.110000 ;
      RECT 1.100000 2232.185000 2225.940000 2233.085000 ;
      RECT 0.000000 2220.540000 2225.940000 2232.185000 ;
      RECT 0.000000 2219.640000 2224.840000 2220.540000 ;
      RECT 0.000000 2178.600000 2225.940000 2219.640000 ;
      RECT 1.100000 2177.700000 2225.940000 2178.600000 ;
      RECT 0.000000 2165.075000 2225.940000 2177.700000 ;
      RECT 0.000000 2164.175000 2224.840000 2165.075000 ;
      RECT 0.000000 2124.210000 2225.940000 2164.175000 ;
      RECT 1.100000 2123.310000 2225.940000 2124.210000 ;
      RECT 0.000000 2109.510000 2225.940000 2123.310000 ;
      RECT 0.000000 2108.610000 2224.840000 2109.510000 ;
      RECT 0.000000 2069.720000 2225.940000 2108.610000 ;
      RECT 1.100000 2068.820000 2225.940000 2069.720000 ;
      RECT 0.000000 2054.040000 2225.940000 2068.820000 ;
      RECT 0.000000 2053.140000 2224.840000 2054.040000 ;
      RECT 0.000000 2015.230000 2225.940000 2053.140000 ;
      RECT 1.100000 2014.330000 2225.940000 2015.230000 ;
      RECT 0.000000 1998.475000 2225.940000 2014.330000 ;
      RECT 0.000000 1997.575000 2224.840000 1998.475000 ;
      RECT 0.000000 1960.840000 2225.940000 1997.575000 ;
      RECT 1.100000 1959.940000 2225.940000 1960.840000 ;
      RECT 0.000000 1943.005000 2225.940000 1959.940000 ;
      RECT 0.000000 1942.105000 2224.840000 1943.005000 ;
      RECT 0.000000 1906.355000 2225.940000 1942.105000 ;
      RECT 1.100000 1905.455000 2225.940000 1906.355000 ;
      RECT 0.000000 1887.540000 2225.940000 1905.455000 ;
      RECT 0.000000 1886.640000 2224.840000 1887.540000 ;
      RECT 0.000000 1851.865000 2225.940000 1886.640000 ;
      RECT 1.100000 1850.965000 2225.940000 1851.865000 ;
      RECT 0.000000 1831.970000 2225.940000 1850.965000 ;
      RECT 0.000000 1831.070000 2224.840000 1831.970000 ;
      RECT 0.000000 1797.475000 2225.940000 1831.070000 ;
      RECT 1.100000 1796.575000 2225.940000 1797.475000 ;
      RECT 0.000000 1776.505000 2225.940000 1796.575000 ;
      RECT 0.000000 1775.605000 2224.840000 1776.505000 ;
      RECT 0.000000 1742.990000 2225.940000 1775.605000 ;
      RECT 1.100000 1742.090000 2225.940000 1742.990000 ;
      RECT 0.000000 1721.035000 2225.940000 1742.090000 ;
      RECT 0.000000 1720.135000 2224.840000 1721.035000 ;
      RECT 0.000000 1688.500000 2225.940000 1720.135000 ;
      RECT 1.100000 1687.600000 2225.940000 1688.500000 ;
      RECT 0.000000 1665.470000 2225.940000 1687.600000 ;
      RECT 0.000000 1664.570000 2224.840000 1665.470000 ;
      RECT 0.000000 1634.110000 2225.940000 1664.570000 ;
      RECT 1.100000 1633.210000 2225.940000 1634.110000 ;
      RECT 0.000000 1610.000000 2225.940000 1633.210000 ;
      RECT 0.000000 1609.100000 2224.840000 1610.000000 ;
      RECT 0.000000 1579.620000 2225.940000 1609.100000 ;
      RECT 1.100000 1578.720000 2225.940000 1579.620000 ;
      RECT 0.000000 1554.535000 2225.940000 1578.720000 ;
      RECT 0.000000 1553.635000 2224.840000 1554.535000 ;
      RECT 0.000000 1525.135000 2225.940000 1553.635000 ;
      RECT 1.100000 1524.235000 2225.940000 1525.135000 ;
      RECT 0.000000 1498.970000 2225.940000 1524.235000 ;
      RECT 0.000000 1498.070000 2224.840000 1498.970000 ;
      RECT 0.000000 1470.745000 2225.940000 1498.070000 ;
      RECT 1.100000 1469.845000 2225.940000 1470.745000 ;
      RECT 0.000000 1443.500000 2225.940000 1469.845000 ;
      RECT 0.000000 1442.600000 2224.840000 1443.500000 ;
      RECT 0.000000 1416.255000 2225.940000 1442.600000 ;
      RECT 1.100000 1415.355000 2225.940000 1416.255000 ;
      RECT 0.000000 1388.030000 2225.940000 1415.355000 ;
      RECT 0.000000 1387.130000 2224.840000 1388.030000 ;
      RECT 0.000000 1361.770000 2225.940000 1387.130000 ;
      RECT 1.100000 1360.870000 2225.940000 1361.770000 ;
      RECT 0.000000 1332.465000 2225.940000 1360.870000 ;
      RECT 0.000000 1331.565000 2224.840000 1332.465000 ;
      RECT 0.000000 1307.380000 2225.940000 1331.565000 ;
      RECT 1.100000 1306.480000 2225.940000 1307.380000 ;
      RECT 0.000000 1277.000000 2225.940000 1306.480000 ;
      RECT 0.000000 1276.100000 2224.840000 1277.000000 ;
      RECT 0.000000 1252.890000 2225.940000 1276.100000 ;
      RECT 1.100000 1251.990000 2225.940000 1252.890000 ;
      RECT 0.000000 1221.430000 2225.940000 1251.990000 ;
      RECT 0.000000 1220.530000 2224.840000 1221.430000 ;
      RECT 0.000000 1198.400000 2225.940000 1220.530000 ;
      RECT 1.100000 1197.500000 2225.940000 1198.400000 ;
      RECT 0.000000 1165.965000 2225.940000 1197.500000 ;
      RECT 0.000000 1165.065000 2224.840000 1165.965000 ;
      RECT 0.000000 1144.010000 2225.940000 1165.065000 ;
      RECT 1.100000 1143.110000 2225.940000 1144.010000 ;
      RECT 0.000000 1110.495000 2225.940000 1143.110000 ;
      RECT 0.000000 1109.595000 2224.840000 1110.495000 ;
      RECT 0.000000 1089.525000 2225.940000 1109.595000 ;
      RECT 1.100000 1088.625000 2225.940000 1089.525000 ;
      RECT 0.000000 1054.930000 2225.940000 1088.625000 ;
      RECT 0.000000 1054.030000 2224.840000 1054.930000 ;
      RECT 0.000000 1035.035000 2225.940000 1054.030000 ;
      RECT 1.100000 1034.135000 2225.940000 1035.035000 ;
      RECT 0.000000 999.460000 2225.940000 1034.135000 ;
      RECT 0.000000 998.560000 2224.840000 999.460000 ;
      RECT 0.000000 980.645000 2225.940000 998.560000 ;
      RECT 1.100000 979.745000 2225.940000 980.645000 ;
      RECT 0.000000 943.995000 2225.940000 979.745000 ;
      RECT 0.000000 943.095000 2224.840000 943.995000 ;
      RECT 0.000000 926.160000 2225.940000 943.095000 ;
      RECT 1.100000 925.260000 2225.940000 926.160000 ;
      RECT 0.000000 888.430000 2225.940000 925.260000 ;
      RECT 0.000000 887.530000 2224.840000 888.430000 ;
      RECT 0.000000 871.670000 2225.940000 887.530000 ;
      RECT 1.100000 870.770000 2225.940000 871.670000 ;
      RECT 0.000000 832.960000 2225.940000 870.770000 ;
      RECT 0.000000 832.060000 2224.840000 832.960000 ;
      RECT 0.000000 817.280000 2225.940000 832.060000 ;
      RECT 1.100000 816.380000 2225.940000 817.280000 ;
      RECT 0.000000 777.490000 2225.940000 816.380000 ;
      RECT 0.000000 776.590000 2224.840000 777.490000 ;
      RECT 0.000000 762.790000 2225.940000 776.590000 ;
      RECT 1.100000 761.890000 2225.940000 762.790000 ;
      RECT 0.000000 721.925000 2225.940000 761.890000 ;
      RECT 0.000000 721.025000 2224.840000 721.925000 ;
      RECT 0.000000 708.305000 2225.940000 721.025000 ;
      RECT 1.100000 707.405000 2225.940000 708.305000 ;
      RECT 0.000000 666.460000 2225.940000 707.405000 ;
      RECT 0.000000 665.560000 2224.840000 666.460000 ;
      RECT 0.000000 653.915000 2225.940000 665.560000 ;
      RECT 1.100000 653.015000 2225.940000 653.915000 ;
      RECT 0.000000 610.890000 2225.940000 653.015000 ;
      RECT 0.000000 609.990000 2224.840000 610.890000 ;
      RECT 0.000000 599.425000 2225.940000 609.990000 ;
      RECT 1.100000 598.525000 2225.940000 599.425000 ;
      RECT 0.000000 555.425000 2225.940000 598.525000 ;
      RECT 0.000000 554.525000 2224.840000 555.425000 ;
      RECT 0.000000 544.940000 2225.940000 554.525000 ;
      RECT 1.100000 544.040000 2225.940000 544.940000 ;
      RECT 0.000000 499.955000 2225.940000 544.040000 ;
      RECT 0.000000 499.055000 2224.840000 499.955000 ;
      RECT 0.000000 490.550000 2225.940000 499.055000 ;
      RECT 1.100000 489.650000 2225.940000 490.550000 ;
      RECT 0.000000 444.390000 2225.940000 489.650000 ;
      RECT 0.000000 443.490000 2224.840000 444.390000 ;
      RECT 0.000000 436.060000 2225.940000 443.490000 ;
      RECT 1.100000 435.160000 2225.940000 436.060000 ;
      RECT 0.000000 388.920000 2225.940000 435.160000 ;
      RECT 0.000000 388.020000 2224.840000 388.920000 ;
      RECT 0.000000 381.570000 2225.940000 388.020000 ;
      RECT 1.100000 380.670000 2225.940000 381.570000 ;
      RECT 0.000000 333.455000 2225.940000 380.670000 ;
      RECT 0.000000 332.555000 2224.840000 333.455000 ;
      RECT 0.000000 327.180000 2225.940000 332.555000 ;
      RECT 1.100000 326.280000 2225.940000 327.180000 ;
      RECT 0.000000 277.890000 2225.940000 326.280000 ;
      RECT 0.000000 276.990000 2224.840000 277.890000 ;
      RECT 0.000000 272.695000 2225.940000 276.990000 ;
      RECT 1.100000 271.795000 2225.940000 272.695000 ;
      RECT 0.000000 222.420000 2225.940000 271.795000 ;
      RECT 0.000000 221.520000 2224.840000 222.420000 ;
      RECT 0.000000 218.205000 2225.940000 221.520000 ;
      RECT 1.100000 217.305000 2225.940000 218.205000 ;
      RECT 0.000000 166.950000 2225.940000 217.305000 ;
      RECT 0.000000 166.050000 2224.840000 166.950000 ;
      RECT 0.000000 163.815000 2225.940000 166.050000 ;
      RECT 1.100000 162.915000 2225.940000 163.815000 ;
      RECT 0.000000 111.385000 2225.940000 162.915000 ;
      RECT 0.000000 110.485000 2224.840000 111.385000 ;
      RECT 0.000000 109.330000 2225.940000 110.485000 ;
      RECT 1.100000 108.430000 2225.940000 109.330000 ;
      RECT 0.000000 55.920000 2225.940000 108.430000 ;
      RECT 0.000000 55.020000 2224.840000 55.920000 ;
      RECT 0.000000 54.840000 2225.940000 55.020000 ;
      RECT 1.100000 53.940000 2225.940000 54.840000 ;
      RECT 0.000000 18.460000 2225.940000 53.940000 ;
      RECT 2212.560000 13.660000 2225.940000 18.460000 ;
      RECT 0.000000 13.660000 13.380000 18.460000 ;
      RECT 0.000000 12.660000 2225.940000 13.660000 ;
      RECT 2218.360000 7.860000 2225.940000 12.660000 ;
      RECT 0.000000 7.860000 7.580000 12.660000 ;
      RECT 0.000000 2.900000 2225.940000 7.860000 ;
      RECT 0.000000 2.000000 2224.840000 2.900000 ;
      RECT 0.000000 1.725000 2225.940000 2.000000 ;
      RECT 1.100000 0.825000 2225.940000 1.725000 ;
      RECT 0.000000 0.000000 2225.940000 0.825000 ;
    LAYER met4 ;
      RECT 0.000000 2885.540000 2225.940000 2895.100000 ;
      RECT 12.380000 2879.740000 2213.560000 2885.540000 ;
      RECT 2212.560000 13.660000 2213.560000 2879.740000 ;
      RECT 18.180000 13.660000 2207.760000 2879.740000 ;
      RECT 12.380000 13.660000 13.380000 2879.740000 ;
      RECT 2218.360000 7.860000 2225.940000 2885.540000 ;
      RECT 12.380000 7.860000 2213.560000 13.660000 ;
      RECT 0.000000 7.860000 7.580000 2885.540000 ;
      RECT 0.000000 0.000000 2225.940000 7.860000 ;
  END
END rest_top

END LIBRARY
